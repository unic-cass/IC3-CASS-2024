// This is the unpowered netlist.
module wb_RAxM (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_sta_o,
    wbs_stb_i,
    wbs_we_i,
    la_data_in,
    la_data_out,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 output wbs_sta_o;
 input wbs_stb_i;
 input wbs_we_i;
 input [47:0] la_data_in;
 output [31:0] la_data_out;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;

 wire net294;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire \mul_la.P_[0] ;
 wire \mul_la.lob_4.A[0] ;
 wire \mul_la.lob_4.B[0] ;
 wire \mul_la.lob_4.L[0] ;
 wire \mul_la.lob_4.L[10] ;
 wire \mul_la.lob_4.L[11] ;
 wire \mul_la.lob_4.L[12] ;
 wire \mul_la.lob_4.L[13] ;
 wire \mul_la.lob_4.L[14] ;
 wire \mul_la.lob_4.L[15] ;
 wire \mul_la.lob_4.L[1] ;
 wire \mul_la.lob_4.L[2] ;
 wire \mul_la.lob_4.L[3] ;
 wire \mul_la.lob_4.L[4] ;
 wire \mul_la.lob_4.L[5] ;
 wire \mul_la.lob_4.L[6] ;
 wire \mul_la.lob_4.L[7] ;
 wire \mul_la.lob_4.L[8] ;
 wire \mul_la.lob_4.L[9] ;
 wire \mul_la.reg_a0[10] ;
 wire \mul_la.reg_a0[11] ;
 wire \mul_la.reg_a0[12] ;
 wire \mul_la.reg_a0[13] ;
 wire \mul_la.reg_a0[14] ;
 wire \mul_la.reg_a0[15] ;
 wire \mul_la.reg_a0[1] ;
 wire \mul_la.reg_a0[2] ;
 wire \mul_la.reg_a0[3] ;
 wire \mul_la.reg_a0[4] ;
 wire \mul_la.reg_a0[5] ;
 wire \mul_la.reg_a0[6] ;
 wire \mul_la.reg_a0[7] ;
 wire \mul_la.reg_a0[8] ;
 wire \mul_la.reg_a0[9] ;
 wire \mul_la.reg_b0[10] ;
 wire \mul_la.reg_b0[11] ;
 wire \mul_la.reg_b0[12] ;
 wire \mul_la.reg_b0[13] ;
 wire \mul_la.reg_b0[14] ;
 wire \mul_la.reg_b0[15] ;
 wire \mul_la.reg_b0[1] ;
 wire \mul_la.reg_b0[2] ;
 wire \mul_la.reg_b0[3] ;
 wire \mul_la.reg_b0[4] ;
 wire \mul_la.reg_b0[5] ;
 wire \mul_la.reg_b0[6] ;
 wire \mul_la.reg_b0[7] ;
 wire \mul_la.reg_b0[8] ;
 wire \mul_la.reg_b0[9] ;
 wire \mul_la.reg_p[10] ;
 wire \mul_la.reg_p[11] ;
 wire \mul_la.reg_p[12] ;
 wire \mul_la.reg_p[13] ;
 wire \mul_la.reg_p[14] ;
 wire \mul_la.reg_p[15] ;
 wire \mul_la.reg_p[16] ;
 wire \mul_la.reg_p[17] ;
 wire \mul_la.reg_p[18] ;
 wire \mul_la.reg_p[19] ;
 wire \mul_la.reg_p[1] ;
 wire \mul_la.reg_p[20] ;
 wire \mul_la.reg_p[21] ;
 wire \mul_la.reg_p[22] ;
 wire \mul_la.reg_p[23] ;
 wire \mul_la.reg_p[24] ;
 wire \mul_la.reg_p[25] ;
 wire \mul_la.reg_p[26] ;
 wire \mul_la.reg_p[27] ;
 wire \mul_la.reg_p[28] ;
 wire \mul_la.reg_p[29] ;
 wire \mul_la.reg_p[2] ;
 wire \mul_la.reg_p[30] ;
 wire \mul_la.reg_p[31] ;
 wire \mul_la.reg_p[3] ;
 wire \mul_la.reg_p[4] ;
 wire \mul_la.reg_p[5] ;
 wire \mul_la.reg_p[6] ;
 wire \mul_la.reg_p[7] ;
 wire \mul_la.reg_p[8] ;
 wire \mul_la.reg_p[9] ;
 wire \mul_wb.P_[0] ;
 wire \mul_wb.a[0] ;
 wire \mul_wb.a[10] ;
 wire \mul_wb.a[11] ;
 wire \mul_wb.a[12] ;
 wire \mul_wb.a[13] ;
 wire \mul_wb.a[14] ;
 wire \mul_wb.a[15] ;
 wire \mul_wb.a[1] ;
 wire \mul_wb.a[2] ;
 wire \mul_wb.a[3] ;
 wire \mul_wb.a[4] ;
 wire \mul_wb.a[5] ;
 wire \mul_wb.a[6] ;
 wire \mul_wb.a[7] ;
 wire \mul_wb.a[8] ;
 wire \mul_wb.a[9] ;
 wire \mul_wb.b[0] ;
 wire \mul_wb.b[10] ;
 wire \mul_wb.b[11] ;
 wire \mul_wb.b[12] ;
 wire \mul_wb.b[13] ;
 wire \mul_wb.b[14] ;
 wire \mul_wb.b[15] ;
 wire \mul_wb.b[1] ;
 wire \mul_wb.b[2] ;
 wire \mul_wb.b[3] ;
 wire \mul_wb.b[4] ;
 wire \mul_wb.b[5] ;
 wire \mul_wb.b[6] ;
 wire \mul_wb.b[7] ;
 wire \mul_wb.b[8] ;
 wire \mul_wb.b[9] ;
 wire \mul_wb.l[0] ;
 wire \mul_wb.l[10] ;
 wire \mul_wb.l[11] ;
 wire \mul_wb.l[12] ;
 wire \mul_wb.l[13] ;
 wire \mul_wb.l[14] ;
 wire \mul_wb.l[15] ;
 wire \mul_wb.l[1] ;
 wire \mul_wb.l[2] ;
 wire \mul_wb.l[3] ;
 wire \mul_wb.l[4] ;
 wire \mul_wb.l[5] ;
 wire \mul_wb.l[6] ;
 wire \mul_wb.l[7] ;
 wire \mul_wb.l[8] ;
 wire \mul_wb.l[9] ;
 wire \mul_wb.lob_4.A[0] ;
 wire \mul_wb.lob_4.B[0] ;
 wire \mul_wb.lob_4.L[0] ;
 wire \mul_wb.lob_4.L[10] ;
 wire \mul_wb.lob_4.L[11] ;
 wire \mul_wb.lob_4.L[12] ;
 wire \mul_wb.lob_4.L[13] ;
 wire \mul_wb.lob_4.L[14] ;
 wire \mul_wb.lob_4.L[15] ;
 wire \mul_wb.lob_4.L[1] ;
 wire \mul_wb.lob_4.L[2] ;
 wire \mul_wb.lob_4.L[3] ;
 wire \mul_wb.lob_4.L[4] ;
 wire \mul_wb.lob_4.L[5] ;
 wire \mul_wb.lob_4.L[6] ;
 wire \mul_wb.lob_4.L[7] ;
 wire \mul_wb.lob_4.L[8] ;
 wire \mul_wb.lob_4.L[9] ;
 wire \mul_wb.p[0] ;
 wire \mul_wb.p[10] ;
 wire \mul_wb.p[11] ;
 wire \mul_wb.p[12] ;
 wire \mul_wb.p[13] ;
 wire \mul_wb.p[14] ;
 wire \mul_wb.p[15] ;
 wire \mul_wb.p[16] ;
 wire \mul_wb.p[17] ;
 wire \mul_wb.p[18] ;
 wire \mul_wb.p[19] ;
 wire \mul_wb.p[1] ;
 wire \mul_wb.p[20] ;
 wire \mul_wb.p[21] ;
 wire \mul_wb.p[22] ;
 wire \mul_wb.p[23] ;
 wire \mul_wb.p[24] ;
 wire \mul_wb.p[25] ;
 wire \mul_wb.p[26] ;
 wire \mul_wb.p[27] ;
 wire \mul_wb.p[28] ;
 wire \mul_wb.p[29] ;
 wire \mul_wb.p[2] ;
 wire \mul_wb.p[30] ;
 wire \mul_wb.p[31] ;
 wire \mul_wb.p[3] ;
 wire \mul_wb.p[4] ;
 wire \mul_wb.p[5] ;
 wire \mul_wb.p[6] ;
 wire \mul_wb.p[7] ;
 wire \mul_wb.p[8] ;
 wire \mul_wb.p[9] ;
 wire \mul_wb.reg_a0[10] ;
 wire \mul_wb.reg_a0[11] ;
 wire \mul_wb.reg_a0[12] ;
 wire \mul_wb.reg_a0[13] ;
 wire \mul_wb.reg_a0[14] ;
 wire \mul_wb.reg_a0[15] ;
 wire \mul_wb.reg_a0[1] ;
 wire \mul_wb.reg_a0[2] ;
 wire \mul_wb.reg_a0[3] ;
 wire \mul_wb.reg_a0[4] ;
 wire \mul_wb.reg_a0[5] ;
 wire \mul_wb.reg_a0[6] ;
 wire \mul_wb.reg_a0[7] ;
 wire \mul_wb.reg_a0[8] ;
 wire \mul_wb.reg_a0[9] ;
 wire \mul_wb.reg_b0[10] ;
 wire \mul_wb.reg_b0[11] ;
 wire \mul_wb.reg_b0[12] ;
 wire \mul_wb.reg_b0[13] ;
 wire \mul_wb.reg_b0[14] ;
 wire \mul_wb.reg_b0[15] ;
 wire \mul_wb.reg_b0[1] ;
 wire \mul_wb.reg_b0[2] ;
 wire \mul_wb.reg_b0[3] ;
 wire \mul_wb.reg_b0[4] ;
 wire \mul_wb.reg_b0[5] ;
 wire \mul_wb.reg_b0[6] ;
 wire \mul_wb.reg_b0[7] ;
 wire \mul_wb.reg_b0[8] ;
 wire \mul_wb.reg_b0[9] ;
 wire \mul_wb.reg_p[10] ;
 wire \mul_wb.reg_p[11] ;
 wire \mul_wb.reg_p[12] ;
 wire \mul_wb.reg_p[13] ;
 wire \mul_wb.reg_p[14] ;
 wire \mul_wb.reg_p[15] ;
 wire \mul_wb.reg_p[16] ;
 wire \mul_wb.reg_p[17] ;
 wire \mul_wb.reg_p[18] ;
 wire \mul_wb.reg_p[19] ;
 wire \mul_wb.reg_p[1] ;
 wire \mul_wb.reg_p[20] ;
 wire \mul_wb.reg_p[21] ;
 wire \mul_wb.reg_p[22] ;
 wire \mul_wb.reg_p[23] ;
 wire \mul_wb.reg_p[24] ;
 wire \mul_wb.reg_p[25] ;
 wire \mul_wb.reg_p[26] ;
 wire \mul_wb.reg_p[27] ;
 wire \mul_wb.reg_p[28] ;
 wire \mul_wb.reg_p[29] ;
 wire \mul_wb.reg_p[2] ;
 wire \mul_wb.reg_p[30] ;
 wire \mul_wb.reg_p[31] ;
 wire \mul_wb.reg_p[3] ;
 wire \mul_wb.reg_p[4] ;
 wire \mul_wb.reg_p[5] ;
 wire \mul_wb.reg_p[6] ;
 wire \mul_wb.reg_p[7] ;
 wire \mul_wb.reg_p[8] ;
 wire \mul_wb.reg_p[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_3325_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(wbs_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(wbs_dat_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(la_data_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(la_data_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(la_data_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(wbs_adr_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(wbs_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(la_data_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A (.DIODE(\mul_wb.lob_4.L[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A (.DIODE(\mul_wb.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A (.DIODE(\mul_wb.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A (.DIODE(\mul_la.lob_4.L[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__D (.DIODE(_3397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__A (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__A (.DIODE(\mul_wb.lob_4.L[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__A (.DIODE(\mul_wb.lob_4.L[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__A1 (.DIODE(\mul_wb.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__B1 (.DIODE(\mul_wb.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__B (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__D (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__D (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__A (.DIODE(\mul_wb.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__A (.DIODE(\mul_wb.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__D (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__B (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__B (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__B (.DIODE(\mul_wb.lob_4.L[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__B (.DIODE(\mul_wb.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__C_N (.DIODE(\mul_wb.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__A (.DIODE(\mul_wb.lob_4.L[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__C_N (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__A1 (.DIODE(\mul_wb.lob_4.L[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A (.DIODE(\mul_wb.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__C (.DIODE(\mul_wb.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__A (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__B (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__A1 (.DIODE(\mul_wb.lob_4.L[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__B2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__C (.DIODE(\mul_wb.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__B2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__A1 (.DIODE(\mul_wb.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__A1 (.DIODE(\mul_wb.lob_4.L[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__B (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__C (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__D (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__C (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A_N (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__C (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__A (.DIODE(\mul_wb.lob_4.L[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__A1 (.DIODE(\mul_wb.lob_4.L[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__B2 (.DIODE(\mul_wb.lob_4.L[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__B (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__A (.DIODE(\mul_wb.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__B (.DIODE(_3397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__C (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__B2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__A (.DIODE(\mul_wb.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__B2 (.DIODE(\mul_wb.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__A1 (.DIODE(\mul_wb.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__B2 (.DIODE(\mul_wb.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__C (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__B1 (.DIODE(\mul_wb.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__A (.DIODE(\mul_wb.lob_4.L[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__A (.DIODE(\mul_wb.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__A1 (.DIODE(\mul_wb.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__A1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__A1 (.DIODE(\mul_wb.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__B1 (.DIODE(\mul_wb.lob_4.L[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__A1 (.DIODE(\mul_wb.lob_4.L[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__B2 (.DIODE(\mul_wb.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__A (.DIODE(_3608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__B (.DIODE(_3613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__B1 (.DIODE(_3614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__C (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__D (.DIODE(_3614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__A (.DIODE(\mul_wb.reg_a0[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__B (.DIODE(_3614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__B2 (.DIODE(\mul_wb.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__B2 (.DIODE(\mul_wb.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__A (.DIODE(\mul_wb.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__D_N (.DIODE(\mul_wb.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__A1 (.DIODE(\mul_wb.lob_4.L[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__B2 (.DIODE(\mul_wb.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__A (.DIODE(\mul_wb.lob_4.L[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__A (.DIODE(\mul_wb.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__A1 (.DIODE(\mul_wb.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__B2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__A (.DIODE(\mul_wb.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__A1 (.DIODE(\mul_wb.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__B1 (.DIODE(\mul_wb.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__B2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A1 (.DIODE(\mul_wb.lob_4.L[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__A (.DIODE(\mul_wb.lob_4.L[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__B (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__B (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__A (.DIODE(\mul_wb.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__A (.DIODE(\mul_wb.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__A1 (.DIODE(\mul_wb.lob_4.L[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__B2 (.DIODE(\mul_wb.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__A (.DIODE(\mul_wb.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__A (.DIODE(_3614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__B (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__B2 (.DIODE(\mul_wb.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__A (.DIODE(\mul_wb.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__B2 (.DIODE(\mul_wb.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__A1 (.DIODE(\mul_wb.lob_4.L[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__B2 (.DIODE(\mul_wb.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__A1 (.DIODE(\mul_wb.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4140__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4140__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__A (.DIODE(\mul_wb.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4146__A (.DIODE(\mul_wb.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__A (.DIODE(\mul_wb.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__A (.DIODE(\mul_wb.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__A (.DIODE(\mul_wb.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A1 (.DIODE(\mul_wb.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__B2 (.DIODE(\mul_wb.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__B2 (.DIODE(\mul_wb.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__A (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__B (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__C_N (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__A1 (.DIODE(_3608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__A2 (.DIODE(_3613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__A (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__A (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__B2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__A (.DIODE(\mul_wb.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__A (.DIODE(\mul_wb.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__C (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__A1 (.DIODE(\mul_wb.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__B2 (.DIODE(\mul_wb.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__B2 (.DIODE(\mul_wb.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__A1 (.DIODE(\mul_wb.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__B2 (.DIODE(\mul_wb.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__A1 (.DIODE(\mul_wb.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__B2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4219__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__C_N (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__A1 (.DIODE(_3608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__A2 (.DIODE(_3613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__B1 (.DIODE(\mul_wb.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__A1 (.DIODE(\mul_wb.lob_4.L[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__B2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__A (.DIODE(\mul_wb.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__A1 (.DIODE(\mul_wb.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__B (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4262__A (.DIODE(\mul_wb.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__B2 (.DIODE(\mul_wb.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__B1 (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__D (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__B1 (.DIODE(\mul_wb.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__A1 (.DIODE(_3614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__C_N (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__A1 (.DIODE(_3608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__A2 (.DIODE(_3613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__A (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4310__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4310__B (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__B1 (.DIODE(\mul_wb.lob_4.L[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__A1 (.DIODE(\mul_wb.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__A1 (.DIODE(\mul_wb.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__B2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__C (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__A1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__B2 (.DIODE(\mul_wb.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__A1 (.DIODE(\mul_wb.lob_4.L[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__A1 (.DIODE(\mul_wb.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__B2 (.DIODE(\mul_wb.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__A1 (.DIODE(\mul_wb.lob_4.L[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__B1 (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__A1 (.DIODE(_3614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__A_N (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__B (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__C (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__A1 (.DIODE(_3608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__A2 (.DIODE(_3613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__C (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__D (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__B2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__B2 (.DIODE(\mul_wb.lob_4.L[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__A (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__A1 (.DIODE(\mul_wb.lob_4.L[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__B2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__B2 (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__A (.DIODE(\mul_wb.lob_4.L[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4384__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__B2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__D (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__A_N (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__B (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__C (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__A (.DIODE(_3614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__A1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__B2 (.DIODE(\mul_wb.lob_4.L[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__B2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__B2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__B (.DIODE(_3683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__C (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__D (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__C_N (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__B2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__D (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__A1 (.DIODE(\mul_wb.lob_4.L[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__B2 (.DIODE(\mul_wb.lob_4.L[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__B2 (.DIODE(_3683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__A (.DIODE(_3683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__C (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__D (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__C_N (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__A (.DIODE(_3657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__A1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__B2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__A (.DIODE(\mul_wb.lob_4.L[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__B1 (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__D (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__A (.DIODE(_3657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__B2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__C (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__D (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__C_N (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__B2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__C (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__D (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__A1 (.DIODE(\mul_wb.lob_4.L[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__B1 (.DIODE(\mul_wb.lob_4.L[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__A (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__A (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__B (.DIODE(_3657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__C (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__D (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__A1 (.DIODE(_3657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__B2 (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__A (.DIODE(_3683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__B2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__B (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__C (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__D (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__C_N (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__A2 (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__B (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__B2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__C (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__D (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__B1 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__A (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__A1 (.DIODE(_3683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__B2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__A (.DIODE(_3587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__B (.DIODE(_3683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__C (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__D (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__B2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__A (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__B2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__C (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__D (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__A2 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__B1 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__C_N (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__A (.DIODE(_3657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__B2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__C (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__D (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__B2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__C (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__B (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__A1 (.DIODE(_3722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__B2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__B (.DIODE(_3722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__C (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__D (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__A (.DIODE(_3587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__B2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__C (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__D (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__A (.DIODE(_3614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__A (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__B (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__C (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__B (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__B1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__A_N (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__A (.DIODE(_0852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__A_N (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__B (.DIODE(_0852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__A2 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__B2 (.DIODE(_3683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__C (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__D (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__B2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__C (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__D (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__B (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__A (.DIODE(_3614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__A (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__B (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__C (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__A1_N (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__A2_N (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__B1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__B (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__B (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__A2 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__A1 (.DIODE(_3587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__A2 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__A (.DIODE(_3722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__B (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__B2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__C (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__D (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__A (.DIODE(_0346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__B (.DIODE(_0442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__B1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__B2 (.DIODE(_3614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__A (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__B (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__C (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__B1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__B (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__B (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__A (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__A (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A1 (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__B1 (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__A2 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A1_N (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A2_N (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A1 (.DIODE(_0346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__B2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__B (.DIODE(_0346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__C (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__D (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__A (.DIODE(_3722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__A2 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__B1 (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__B2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__C (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__D (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__B (.DIODE(_0442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__B (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__A1 (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__A2 (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__B1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__A2 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__B1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__B2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__C (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__D (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__B (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A2 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__B2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__C (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__D (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__B (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__B2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__C (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__D (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A (.DIODE(_0442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A2 (.DIODE(_0442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__B1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__B1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__C1 (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A1_N (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A1 (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A3 (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__B1 (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__A (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__C (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__D (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__A1_N (.DIODE(_3722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__A2_N (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__B2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__A (.DIODE(_0346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__C (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__D (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__B (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__B (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__B (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__B1 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__B (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__A2 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__B (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__A2 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A2 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__B2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__C (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__D (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A (.DIODE(_0346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__B2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__C (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__D (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__B (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__B1 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__A2_N (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A1 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__B (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A2 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__B1 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__C1 (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__B (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__B1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__B2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__B2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__C (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__D (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__A1 (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__B1 (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__B1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__B2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__C (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__D (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__A2 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__B (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__B1 (.DIODE(_0346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__B2 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__B (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__C (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__D_N (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A1 (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__A1 (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__A2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__C (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__D (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A (.DIODE(_0442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A1 (.DIODE(_0442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__B1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__B2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__C (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__D (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A2_N (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A2 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__B (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__B (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__C (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__D (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A1 (.DIODE(_0442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A2 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__B1 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__B2 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__C (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__D (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__B (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__A1 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__A (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__B (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__A2 (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__A (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__C_N (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A2_N (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__B1 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__B (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__B1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A3 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A2 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__B1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__B2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__C (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__D (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__A2 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A2 (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__B2 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__B (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__B1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__B2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__A2 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__A_N (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__C (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__A (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__B (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__A2 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A2 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__B1 (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__A1 (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__A2 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__B1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__B1 (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__B1 (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A2 (.DIODE(_3397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__B1_N (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A (.DIODE(\mul_la.lob_4.L[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A (.DIODE(\mul_la.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A (.DIODE(\mul_la.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__A (.DIODE(\mul_la.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__C1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__A (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A (.DIODE(\mul_la.lob_4.L[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__A (.DIODE(\mul_la.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__C (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__B (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__D (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A (.DIODE(\mul_la.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A2 (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__B (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__B1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__B (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__C (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__A (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A (.DIODE(\mul_la.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__B (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__A1 (.DIODE(\mul_la.lob_4.L[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__A2 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__B2 (.DIODE(\mul_la.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__A (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A2 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__B2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A_N (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__A_N (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__C (.DIODE(\mul_la.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__B2 (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A_N (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__B (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A_N (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__A1 (.DIODE(\mul_la.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__B2 (.DIODE(\mul_la.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__A1 (.DIODE(\mul_la.lob_4.L[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A2 (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__B2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A2 (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__B2 (.DIODE(\mul_la.lob_4.L[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A_N (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__B (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A1 (.DIODE(\mul_la.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__A1 (.DIODE(\mul_la.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A2 (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__B1 (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A2 (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__B1 (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A (.DIODE(\mul_la.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A (.DIODE(\mul_la.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__B2 (.DIODE(\mul_la.lob_4.L[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A1 (.DIODE(\mul_la.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__B1 (.DIODE(\mul_la.lob_4.L[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__A1 (.DIODE(\mul_la.lob_4.L[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__B (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__A1 (.DIODE(\mul_la.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__A (.DIODE(_1794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__B (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__A (.DIODE(_1794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__B (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__B2 (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__B (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__C (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__A (.DIODE(\mul_la.reg_a0[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__B1 (.DIODE(\mul_la.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__A (.DIODE(\mul_la.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__A1 (.DIODE(\mul_la.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__B2 (.DIODE(\mul_la.lob_4.L[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__A1 (.DIODE(\mul_la.lob_4.L[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__B2 (.DIODE(\mul_la.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__C (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__B2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__A (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__B (.DIODE(_1829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__A (.DIODE(\mul_la.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__A2 (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__A1 (.DIODE(\mul_la.lob_4.L[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__B2 (.DIODE(\mul_la.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__A1 (.DIODE(\mul_la.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__A2 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__B2 (.DIODE(\mul_la.lob_4.L[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__B2 (.DIODE(\mul_la.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__B (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__B1 (.DIODE(\mul_la.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__A (.DIODE(\mul_la.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A (.DIODE(\mul_la.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__A1 (.DIODE(\mul_la.lob_4.L[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__B2 (.DIODE(\mul_la.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5877__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5879__A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A (.DIODE(\mul_la.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A1 (.DIODE(\mul_la.lob_4.L[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__B1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__A1 (.DIODE(\mul_la.lob_4.L[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__B1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__A (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__A (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__B (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__B (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__B2 (.DIODE(\mul_la.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__A1 (.DIODE(\mul_la.lob_4.L[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__A2 (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__B2 (.DIODE(\mul_la.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__B (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A1 (.DIODE(\mul_la.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__B2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__A1 (.DIODE(\mul_la.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__B2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__A2_N (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__B1 (.DIODE(_1890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__A_N (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__B (.DIODE(_1890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__A (.DIODE(\mul_la.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__A1 (.DIODE(\mul_la.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__B2 (.DIODE(\mul_la.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__B2 (.DIODE(\mul_la.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__A_N (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__C (.DIODE(_1876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__D (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A2 (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__B1 (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__B2 (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__A (.DIODE(_1829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__A (.DIODE(\mul_la.lob_4.L[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__A (.DIODE(\mul_la.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__A1 (.DIODE(\mul_la.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__B (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__B2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__A1 (.DIODE(\mul_la.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__A2 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__A2 (.DIODE(_1890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__B1 (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__C (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__D (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__A2 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__A1_N (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__A1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__A2 (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__B1 (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__C1 (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__B (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__A1 (.DIODE(\mul_la.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__B2 (.DIODE(\mul_la.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__B2 (.DIODE(\mul_la.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__A (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__A (.DIODE(_1829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__B (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__A2 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__B2 (.DIODE(\mul_la.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__B1 (.DIODE(\mul_la.lob_4.L[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__B2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__A1 (.DIODE(\mul_la.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__B (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__B2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__A1 (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__A2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__B1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__A1 (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__A2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__B1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__A2 (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__B1 (.DIODE(_1978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__C (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__D (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__A1 (.DIODE(\mul_la.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__B2 (.DIODE(\mul_la.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__A (.DIODE(\mul_la.lob_4.L[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__A1 (.DIODE(\mul_la.lob_4.L[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__A (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__B (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6027__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6027__B (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__A (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__B (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__B (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A (.DIODE(_1829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__B2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__B (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__C (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__A (.DIODE(\mul_la.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__A1 (.DIODE(\mul_la.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__B2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__A1 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__A2 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__B1 (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__A1 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__A2 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__B1 (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__A2 (.DIODE(_1978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__B1 (.DIODE(_2024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__C (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__D (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__A (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__B2 (.DIODE(\mul_la.lob_4.L[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__A1 (.DIODE(\mul_la.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__B2 (.DIODE(\mul_la.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__A (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__B (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__B (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__A2 (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__B (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__A1 (.DIODE(_1890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__B1 (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__B2 (.DIODE(_1876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__A (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__B (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__C (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__D (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__A (.DIODE(_1829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__B (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__A1 (.DIODE(\mul_la.lob_4.L[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__B1 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__B2 (.DIODE(\mul_la.lob_4.L[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__B (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__C (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__A2 (.DIODE(_2024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__B1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__C (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__D_N (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__B2 (.DIODE(\mul_la.lob_4.L[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__A1 (.DIODE(\mul_la.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__B2 (.DIODE(\mul_la.lob_4.L[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__A (.DIODE(_2115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__A (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A2 (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__B1 (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__C1 (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__B (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__A (.DIODE(_1890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__B (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__A2 (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__B1 (.DIODE(_1978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__B2 (.DIODE(_1876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__A (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__B (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__C (.DIODE(_1934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__D (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__B (.DIODE(_2024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__A1 (.DIODE(_1794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__A2 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__B (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__B (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A_N (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__C (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__B (.DIODE(_2141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__C (.DIODE(_2141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__B1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__A1 (.DIODE(\mul_la.lob_4.L[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__B2 (.DIODE(\mul_la.lob_4.L[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__A (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__B (.DIODE(_2176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__A2 (.DIODE(_2061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__B (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A (.DIODE(_1890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__B (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__B (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__A2 (.DIODE(_1978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__B1 (.DIODE(_2024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__B2 (.DIODE(_1876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__A (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__B (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__C (.DIODE(_1979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__D (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A1 (.DIODE(_1794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A2 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__B1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__A2 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__B2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__B2 (.DIODE(\mul_la.lob_4.L[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__B2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__B1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__B1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__B (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6227__C (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__A2 (.DIODE(_2024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__B (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__A1 (.DIODE(\mul_la.lob_4.L[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__B2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__6257__A (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6257__B (.DIODE(_2235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__A2 (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__A (.DIODE(_1890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__B (.DIODE(_2061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6266__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6266__B (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__A2 (.DIODE(_2024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__B2 (.DIODE(_1876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__A (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__B (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__C (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__D_N (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__B (.DIODE(_2141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6280__A1 (.DIODE(_1794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6280__A2 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6280__B1 (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6281__B (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6282__A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__B (.DIODE(_2264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__C (.DIODE(_2264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6291__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6291__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__A (.DIODE(_1809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6319__B1 (.DIODE(_1809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__A (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__B (.DIODE(_2176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__A2 (.DIODE(_2234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__A2 (.DIODE(_2234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__B (.DIODE(_2234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A1 (.DIODE(_1890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A2 (.DIODE(_2061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__A (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__B (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__B (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__B (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__A (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__A (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6355__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6355__B (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__A1 (.DIODE(_1794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__A2 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__B1 (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__B1 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__B1 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__C (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__A2 (.DIODE(_2141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__A (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__B (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__A1 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__A2 (.DIODE(_2176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__B1 (.DIODE(_2235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__A_N (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__B (.DIODE(_1890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__C (.DIODE(_2175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__D (.DIODE(_2234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__A1 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6415__A1 (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6415__A2 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6415__B1 (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6415__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__B (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__C (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__D (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__A (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__B (.DIODE(_2141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__A (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__C (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__A (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__B (.DIODE(_2141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__C (.DIODE(_2401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__B (.DIODE(_2401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__A (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__A1 (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__B (.DIODE(_2264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__A1 (.DIODE(_1794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__A2 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__B1 (.DIODE(_2339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__B (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__C (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__A2 (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__A1 (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__A2 (.DIODE(_2376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6472__B2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__A (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__C (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__D (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__A2 (.DIODE(_2376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__B1 (.DIODE(_2449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__B2 (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__A1 (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__A2 (.DIODE(_2175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__B1 (.DIODE(_2234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__B2 (.DIODE(_1890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__A (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__C (.DIODE(_2176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__D (.DIODE(_2235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__A2 (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__A2 (.DIODE(_2115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__A1 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__A2 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__B1 (.DIODE(_2061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__C1 (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6494__A (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__A (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__B (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__B (.DIODE(_2115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__A2 (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__B1 (.DIODE(_2264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__B2 (.DIODE(_1876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__A (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__B (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__C (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__D (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__A1 (.DIODE(_1794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__A2 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__B1 (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__B (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__C (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__A2 (.DIODE(_2264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6544__A1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6544__A2 (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6544__B1 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6544__C1 (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6545__A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6545__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6548__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6549__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__A (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__B1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__6553__A1 (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6553__A2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6553__B1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6553__C1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__A (.DIODE(_2527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6555__A (.DIODE(_2527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__A (.DIODE(_2527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__A (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__A2 (.DIODE(_2115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__A1_N (.DIODE(_2061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__B1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__B2 (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__A (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__B (.DIODE(_2061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__D (.DIODE(_2141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__A (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__B (.DIODE(_2115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6573__B1 (.DIODE(_2024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__A2 (.DIODE(_2264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__B1 (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__B2 (.DIODE(_1876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__A (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__B (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__C (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__D (.DIODE(_2339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__B (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__B (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__A1 (.DIODE(_1794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__A2 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__B1 (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__B (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__B (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__C (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__A2 (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__A (.DIODE(_1809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__B1 (.DIODE(_1809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__A1 (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__A2 (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__A1 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__B1 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__A_N (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__B (.DIODE(_1890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__C (.DIODE(_2376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__D (.DIODE(_2449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A1 (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__B1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__C1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__A1 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__A2 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__B1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__C1 (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__B (.DIODE(_2303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__A1 (.DIODE(_2061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__A2 (.DIODE(_2141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__B1 (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__B2 (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__A (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__B (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__C (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__D (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__A (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__B (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__B (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__B (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__B (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__B (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__A2 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__B1 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__A2 (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__A2 (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__A1 (.DIODE(_1934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__B1 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__B2 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__A (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__B (.DIODE(_1934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__C (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__D (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__A1 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__A2 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__B1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__C1 (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__B (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__A (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__B (.DIODE(_2235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__A1 (.DIODE(_2061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__A2 (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__B1 (.DIODE(_2264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__B2 (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__A (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__B (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__C (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__D (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__A3 (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__B1 (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__B1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__C1 (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__D1 (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__A (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__A2 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__B1 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__A (.DIODE(_1809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__A2 (.DIODE(_2524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__A2 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__A1 (.DIODE(_1978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__A2 (.DIODE(_2376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__B1 (.DIODE(_2449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__B2 (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__C (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__D (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__A (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__A1 (.DIODE(_2141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__B1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__B (.DIODE(_2141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__C (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__D (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__B (.DIODE(_2141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__C (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__D (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__A (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__C (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6789__A1 (.DIODE(_2024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6789__A2 (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__A1 (.DIODE(_2061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__A2 (.DIODE(_2264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__B1 (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__B2 (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__A (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__B (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__C (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__D (.DIODE(_2339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__B (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__A3 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__B1 (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__B1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__C1 (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__D1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__A (.DIODE(_1877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__B (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__C (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__B (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__B2 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6842__B1 (.DIODE(_1809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__A1 (.DIODE(_1890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__A2 (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__A1 (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__A2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__B1 (.DIODE(_2449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__C1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__A1 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__A2 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__B1 (.DIODE(_2376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__C1 (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__B1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__B1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__B (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__A1 (.DIODE(_2024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__A2 (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__A3 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__B1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__B (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__A1 (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__A2 (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__A1 (.DIODE(_2061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__A2 (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__B1 (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__B2 (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__A (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__B (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__C (.DIODE(_2339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__D (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__B (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__B1 (.DIODE(_1809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6912__B1 (.DIODE(_1809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6917__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6917__B2 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__A1 (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__A2 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__B1 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6920__B1 (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__B1 (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__B (.DIODE(_2339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__A1 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__A2 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__B1 (.DIODE(_2449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__C1 (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__B (.DIODE(_2376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__A (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__B (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6941__B1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__6941__C1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6942__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6971__A1 (.DIODE(_2061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6971__A2 (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__A1 (.DIODE(_2061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__A2 (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__B1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__B2 (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__A (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__B (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__C (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6975__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6975__B (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6976__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6976__B (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__B (.DIODE(_2449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6986__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6987__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6987__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__A (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6992__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__6993__B1 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6993__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6996__A (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6996__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6998__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__7008__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__7008__A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__7011__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__7011__B2 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7022__A (.DIODE(_2989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7022__B (.DIODE(_2990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7024__A (.DIODE(_2989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7024__B (.DIODE(_2990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7034__A (.DIODE(_1809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7036__A1 (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7036__B2 (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7037__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__7037__B (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__A2 (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__A1 (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__A2 (.DIODE(_2376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__B1 (.DIODE(_2449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__B2 (.DIODE(_2141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__B (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__C (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__D (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7047__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__B1 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__B (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__A (.DIODE(_2235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__B (.DIODE(_2339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7053__A (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7053__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__7055__A1 (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7055__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__7071__A1 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7071__A2 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__A (.DIODE(_3047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7082__A (.DIODE(_3047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7082__B (.DIODE(_3049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7086__B1 (.DIODE(_1809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__A2 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__B1 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__B2 (.DIODE(_2061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7091__A1 (.DIODE(_2264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7091__A2 (.DIODE(_2376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7091__B1 (.DIODE(_2449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7091__B2 (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7092__A (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7092__B (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7092__D (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7094__A (.DIODE(_2141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7096__A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__7096__A2 (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7096__B1 (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7096__B2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__C (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__D (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__A (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7101__A1 (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7101__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__B1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__B2 (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__B1 (.DIODE(_3049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7132__B1 (.DIODE(_1809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__B1 (.DIODE(_1809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7137__A1 (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7137__A2 (.DIODE(_2376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7137__B1 (.DIODE(_2449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7137__B2 (.DIODE(_2264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7138__A (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7138__B (.DIODE(_2339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7138__D (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7140__A (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7140__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__7142__A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__7142__A2 (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7142__B1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7142__B2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__7143__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__7143__B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__7143__C (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7143__D (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7145__A (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7145__B (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7156__B1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__7160__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__7160__A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__7163__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__7163__A2 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7175__A1 (.DIODE(_2376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7175__A2 (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7175__B1 (.DIODE(_2449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7175__B2 (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7176__A (.DIODE(_2339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7176__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__7176__C (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7176__D (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7178__A (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7178__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__7180__A1 (.DIODE(_2235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7180__B2 (.DIODE(_2176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7181__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__7181__B (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7182__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__7182__A2 (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7194__A1 (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7194__A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__7197__A (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7197__B (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7219__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__7221__A1 (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7221__A2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7221__B1 (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7221__B2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__7222__A (.DIODE(_2376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7222__B (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7222__C (.DIODE(_2449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7222__D (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7224__A (.DIODE(_2339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7224__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__A1 (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__A2 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__B1 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__B2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__7237__A (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7237__B (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7250__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__7252__A1 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7252__A2 (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7252__B2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__7253__A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__7253__B (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7253__C (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7255__A (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7255__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__7257__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__7265__B1 (.DIODE(_2339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7265__B2 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7285__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__7291__A (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7291__B (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7292__A1 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7292__B2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__7293__A1 (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7293__A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__7294__C (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7311__B1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__7312__A (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7313__B (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7314__A1 (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7314__A2 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7314__B2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7325__A (.DIODE(_3285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7326__D (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7327__B1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__7328__A (.DIODE(_3285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7329__A1 (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7329__A2 (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7329__B1 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7332__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__7333__A (.DIODE(_3291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7334__C (.DIODE(_3285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7335__C_N (.DIODE(_3293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7336__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__7336__B (.DIODE(_3294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7337__A3 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7337__B1 (.DIODE(_3294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7337__B2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__7348__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7348__C (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__7349__B (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__7353__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__7354__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7355__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__7356__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7357__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__7358__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7359__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__7360__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7361__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__7362__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__7363__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__7364__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__7365__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__7366__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7367__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__7368__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__7369__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__7370__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__7371__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__7372__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__7373__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__7374__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__7375__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__7376__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__7377__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__7378__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__7379__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__7380__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__7381__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__7382__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__7383__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__7384__A (.DIODE(_0000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7385__B (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__7388__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7389__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__7390__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7391__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7392__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7393__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7394__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7395__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__7396__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7397__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__7398__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7399__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__7400__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7401__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__7402__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7403__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__7404__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7405__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__7406__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7407__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__7408__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7409__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__7410__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7411__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__7412__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7413__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__7414__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7415__A (.DIODE(_0000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7416__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7417__A (.DIODE(_0000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7418__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7419__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__7421__S (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7422__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__7423__S (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7424__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7425__S (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7426__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7427__S (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7428__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7429__S (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7430__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7431__S (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7432__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7433__S (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7434__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7435__S (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7436__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7437__S (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7438__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__7439__S (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7440__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__7441__S (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7442__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__7443__S (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7444__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__7445__S (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7446__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__7447__S (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7448__A (.DIODE(_0000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7449__S (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7450__A (.DIODE(_0000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7451__S (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7452__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__7454__C (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7455__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7455__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7456__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7456__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7457__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7457__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7458__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7458__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7459__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7459__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7460__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7460__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7461__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7461__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7462__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7462__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7463__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7463__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7464__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7464__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7465__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7465__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7466__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7466__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7467__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7467__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7468__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__7468__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__7469__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__7469__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__7470__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__7470__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__7471__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__7471__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__7472__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__7472__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__7473__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__7473__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__7474__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__7474__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__7475__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__7475__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__7476__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__7476__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__7477__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__7477__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__7478__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__7478__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__7479__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__7479__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__7480__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__7480__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__7481__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__7481__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__7482__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__7482__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__7483__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__7483__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__7484__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7484__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7485__A2 (.DIODE(_3361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7485__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7486__A2 (.DIODE(_3361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7486__B1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__7511__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__7512__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__7513__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__7514__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__7515__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__7516__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__7517__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__7519__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__7520__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__7521__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__7523__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__7525__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__7527__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__7531__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__7532__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__7534__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__7535__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__7536__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__7538__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__7546__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__7548__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__7550__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__7551__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__7552__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__7553__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__7554__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__7555__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__7556__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__7557__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__7559__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__7563__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__7564__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__7566__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__7567__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__7568__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__7569__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__7570__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__7571__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__7572__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__7573__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__7574__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__7598__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__7599__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__7600__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__7601__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__7602__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__7603__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__7604__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__7605__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__7606__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__7607__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__7608__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__7609__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__7610__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__7611__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__7612__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__7613__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__7614__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__7615__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__7616__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__7621__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__7622__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__7623__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__7624__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__7625__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__7626__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__7627__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__7628__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__7629__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__7630__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__7631__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__7632__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__7633__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__7634__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__7635__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__7636__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__7637__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__7638__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__7639__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__7640__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__7641__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__7727__RESET_B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7740__D (.DIODE(\mul_wb.reg_p[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(_1979_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(_1934_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(_3657_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(_3587_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(_2303_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(_2115_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(_2085_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(_2085_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(_0442_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(_0346_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(_0332_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(_0332_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(_3783_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(_3783_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(_3722_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(_3683_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(_2234_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(_2175_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(_2524_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(\mul_la.reg_a0[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(\mul_la.lob_4.L[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(\mul_la.lob_4.L[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(\mul_la.lob_4.L[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(\mul_la.lob_4.L[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(\mul_la.lob_4.L[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_A (.DIODE(\mul_wb.reg_a0[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(\mul_wb.lob_4.L[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_A (.DIODE(\mul_wb.lob_4.L[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_A (.DIODE(\mul_wb.lob_4.L[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(_3361_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(_0000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(_0000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout287_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout288_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout289_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout291_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout292_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold104_A (.DIODE(_3362_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold409_A (.DIODE(\mul_wb.reg_a0[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold410_A (.DIODE(\mul_la.reg_a0[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap211_A (.DIODE(_3613_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap247_A (.DIODE(_3397_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire212_A (.DIODE(_3608_));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_84 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _3791_ (.A(\mul_wb.lob_4.A[0] ),
    .Y(_3363_));
 sky130_fd_sc_hd__inv_2 _3792_ (.A(net269),
    .Y(_3364_));
 sky130_fd_sc_hd__inv_2 _3793_ (.A(net270),
    .Y(_3365_));
 sky130_fd_sc_hd__inv_2 _3794_ (.A(net272),
    .Y(_3366_));
 sky130_fd_sc_hd__inv_2 _3795_ (.A(\mul_wb.lob_4.L[12] ),
    .Y(_3367_));
 sky130_fd_sc_hd__inv_2 _3796_ (.A(net274),
    .Y(_3368_));
 sky130_fd_sc_hd__inv_2 _3797_ (.A(net275),
    .Y(_3369_));
 sky130_fd_sc_hd__inv_2 _3798_ (.A(\mul_wb.lob_4.L[9] ),
    .Y(_3370_));
 sky130_fd_sc_hd__inv_2 _3799_ (.A(\mul_wb.lob_4.L[8] ),
    .Y(_3371_));
 sky130_fd_sc_hd__inv_2 _3800_ (.A(net256),
    .Y(_3372_));
 sky130_fd_sc_hd__inv_2 _3801_ (.A(net259),
    .Y(_3373_));
 sky130_fd_sc_hd__inv_2 _3802_ (.A(net261),
    .Y(_3374_));
 sky130_fd_sc_hd__inv_2 _3803_ (.A(\mul_la.lob_4.L[3] ),
    .Y(_3375_));
 sky130_fd_sc_hd__clkinv_4 _3804_ (.A(net707),
    .Y(_3376_));
 sky130_fd_sc_hd__inv_2 _3805_ (.A(net281),
    .Y(_0000_));
 sky130_fd_sc_hd__or4_4 _3806_ (.A(\mul_wb.reg_a0[2] ),
    .B(\mul_wb.reg_a0[1] ),
    .C(\mul_wb.lob_4.A[0] ),
    .D(\mul_wb.reg_a0[3] ),
    .X(_3377_));
 sky130_fd_sc_hd__or4_4 _3807_ (.A(\mul_wb.reg_a0[4] ),
    .B(\mul_wb.reg_a0[5] ),
    .C(\mul_wb.reg_a0[6] ),
    .D(\mul_wb.reg_a0[7] ),
    .X(_3378_));
 sky130_fd_sc_hd__o41a_4 _3808_ (.A1(\mul_wb.reg_a0[8] ),
    .A2(\mul_wb.reg_a0[9] ),
    .A3(_3377_),
    .A4(_3378_),
    .B1(net266),
    .X(_3379_));
 sky130_fd_sc_hd__and2_1 _3809_ (.A(net266),
    .B(\mul_wb.reg_a0[10] ),
    .X(_3380_));
 sky130_fd_sc_hd__o21ai_4 _3810_ (.A1(_3379_),
    .A2(_3380_),
    .B1(\mul_wb.reg_a0[11] ),
    .Y(_3381_));
 sky130_fd_sc_hd__or3_4 _3811_ (.A(\mul_wb.reg_a0[11] ),
    .B(_3379_),
    .C(_3380_),
    .X(_3382_));
 sky130_fd_sc_hd__and2_4 _3812_ (.A(_3381_),
    .B(_3382_),
    .X(_3383_));
 sky130_fd_sc_hd__nand2_2 _3813_ (.A(_3381_),
    .B(_3382_),
    .Y(_3384_));
 sky130_fd_sc_hd__or4_2 _3814_ (.A(\mul_wb.reg_a0[8] ),
    .B(\mul_wb.reg_a0[9] ),
    .C(\mul_wb.reg_a0[10] ),
    .D(\mul_wb.reg_a0[11] ),
    .X(_3385_));
 sky130_fd_sc_hd__o31a_2 _3815_ (.A1(_3377_),
    .A2(_3378_),
    .A3(_3385_),
    .B1(net266),
    .X(_3386_));
 sky130_fd_sc_hd__o41a_4 _3816_ (.A1(\mul_wb.reg_a0[12] ),
    .A2(_3377_),
    .A3(_3378_),
    .A4(_3385_),
    .B1(net266),
    .X(_3387_));
 sky130_fd_sc_hd__xor2_4 _3817_ (.A(\mul_wb.reg_a0[13] ),
    .B(_3387_),
    .X(_3388_));
 sky130_fd_sc_hd__xnor2_4 _3818_ (.A(\mul_wb.reg_a0[13] ),
    .B(_3387_),
    .Y(_3389_));
 sky130_fd_sc_hd__xor2_4 _3819_ (.A(\mul_wb.reg_a0[12] ),
    .B(_3386_),
    .X(_3390_));
 sky130_fd_sc_hd__nor2_1 _3820_ (.A(_3388_),
    .B(_3390_),
    .Y(_3391_));
 sky130_fd_sc_hd__or2_1 _3821_ (.A(net992),
    .B(\mul_wb.reg_a0[13] ),
    .X(_3392_));
 sky130_fd_sc_hd__or4_1 _3822_ (.A(_3377_),
    .B(_3378_),
    .C(_3385_),
    .D(net993),
    .X(_3393_));
 sky130_fd_sc_hd__o41a_2 _3823_ (.A1(_3377_),
    .A2(_3378_),
    .A3(_3385_),
    .A4(_3392_),
    .B1(net266),
    .X(_3394_));
 sky130_fd_sc_hd__xor2_1 _3824_ (.A(\mul_wb.reg_a0[14] ),
    .B(_3394_),
    .X(_3395_));
 sky130_fd_sc_hd__xnor2_4 _3825_ (.A(\mul_wb.reg_a0[14] ),
    .B(_3394_),
    .Y(_3396_));
 sky130_fd_sc_hd__nor3b_4 _3826_ (.A(net706),
    .B(net994),
    .C_N(net266),
    .Y(_3397_));
 sky130_fd_sc_hd__nor2_1 _3827_ (.A(net249),
    .B(net247),
    .Y(_3398_));
 sky130_fd_sc_hd__nor4_4 _3828_ (.A(_3388_),
    .B(net250),
    .C(net248),
    .D(net247),
    .Y(_3399_));
 sky130_fd_sc_hd__or4_4 _3829_ (.A(_3388_),
    .B(net250),
    .C(net248),
    .D(_3397_),
    .X(_3400_));
 sky130_fd_sc_hd__xor2_2 _3830_ (.A(\mul_wb.reg_a0[10] ),
    .B(_3379_),
    .X(_3401_));
 sky130_fd_sc_hd__xnor2_2 _3831_ (.A(\mul_wb.reg_a0[10] ),
    .B(_3379_),
    .Y(_3402_));
 sky130_fd_sc_hd__o21a_2 _3832_ (.A1(_3377_),
    .A2(_3378_),
    .B1(net266),
    .X(_3403_));
 sky130_fd_sc_hd__o31a_2 _3833_ (.A1(\mul_wb.reg_a0[8] ),
    .A2(_3377_),
    .A3(_3378_),
    .B1(net266),
    .X(_3404_));
 sky130_fd_sc_hd__xor2_4 _3834_ (.A(\mul_wb.reg_a0[9] ),
    .B(_3404_),
    .X(_3405_));
 sky130_fd_sc_hd__xnor2_1 _3835_ (.A(\mul_wb.reg_a0[9] ),
    .B(_3404_),
    .Y(_3406_));
 sky130_fd_sc_hd__nor2_2 _3836_ (.A(net246),
    .B(_3405_),
    .Y(_3407_));
 sky130_fd_sc_hd__xor2_4 _3837_ (.A(\mul_wb.reg_a0[8] ),
    .B(_3403_),
    .X(_3408_));
 sky130_fd_sc_hd__xnor2_2 _3838_ (.A(\mul_wb.reg_a0[8] ),
    .B(_3403_),
    .Y(_3409_));
 sky130_fd_sc_hd__a2111oi_2 _3839_ (.A1(_3381_),
    .A2(_3382_),
    .B1(net246),
    .C1(_3405_),
    .D1(_3408_),
    .Y(_3410_));
 sky130_fd_sc_hd__a2111o_2 _3840_ (.A1(_3381_),
    .A2(_3382_),
    .B1(net246),
    .C1(_3405_),
    .D1(_3408_),
    .X(_3411_));
 sky130_fd_sc_hd__nor2_2 _3841_ (.A(_3400_),
    .B(_3411_),
    .Y(_3412_));
 sky130_fd_sc_hd__o31a_2 _3842_ (.A1(\mul_wb.reg_a0[4] ),
    .A2(\mul_wb.reg_a0[5] ),
    .A3(_3377_),
    .B1(net266),
    .X(_3413_));
 sky130_fd_sc_hd__o41a_2 _3843_ (.A1(\mul_wb.reg_a0[4] ),
    .A2(\mul_wb.reg_a0[5] ),
    .A3(\mul_wb.reg_a0[6] ),
    .A4(_3377_),
    .B1(net266),
    .X(_3414_));
 sky130_fd_sc_hd__xor2_4 _3844_ (.A(\mul_wb.reg_a0[7] ),
    .B(_3414_),
    .X(_3415_));
 sky130_fd_sc_hd__inv_2 _3845_ (.A(_3415_),
    .Y(_3416_));
 sky130_fd_sc_hd__xor2_4 _3846_ (.A(\mul_wb.reg_a0[6] ),
    .B(_3413_),
    .X(_3417_));
 sky130_fd_sc_hd__xnor2_2 _3847_ (.A(\mul_wb.reg_a0[6] ),
    .B(_3413_),
    .Y(_3418_));
 sky130_fd_sc_hd__nor2_1 _3848_ (.A(_3415_),
    .B(_3417_),
    .Y(_3419_));
 sky130_fd_sc_hd__o21a_2 _3849_ (.A1(\mul_wb.reg_a0[1] ),
    .A2(\mul_wb.lob_4.A[0] ),
    .B1(net266),
    .X(_3420_));
 sky130_fd_sc_hd__xor2_4 _3850_ (.A(\mul_wb.reg_a0[2] ),
    .B(_3420_),
    .X(_3421_));
 sky130_fd_sc_hd__xnor2_1 _3851_ (.A(\mul_wb.reg_a0[2] ),
    .B(_3420_),
    .Y(_3422_));
 sky130_fd_sc_hd__o31a_2 _3852_ (.A1(\mul_wb.reg_a0[2] ),
    .A2(\mul_wb.reg_a0[1] ),
    .A3(\mul_wb.lob_4.A[0] ),
    .B1(net266),
    .X(_3423_));
 sky130_fd_sc_hd__xor2_4 _3853_ (.A(\mul_wb.reg_a0[3] ),
    .B(_3423_),
    .X(_3424_));
 sky130_fd_sc_hd__xnor2_1 _3854_ (.A(\mul_wb.reg_a0[3] ),
    .B(_3423_),
    .Y(_3425_));
 sky130_fd_sc_hd__o41a_2 _3855_ (.A1(\mul_wb.reg_a0[2] ),
    .A2(\mul_wb.reg_a0[1] ),
    .A3(\mul_wb.lob_4.A[0] ),
    .A4(\mul_wb.reg_a0[3] ),
    .B1(net266),
    .X(_3426_));
 sky130_fd_sc_hd__o211ai_2 _3856_ (.A1(\mul_wb.reg_a0[4] ),
    .A2(_3377_),
    .B1(\mul_wb.reg_a0[5] ),
    .C1(net266),
    .Y(_3427_));
 sky130_fd_sc_hd__a211o_1 _3857_ (.A1(net266),
    .A2(\mul_wb.reg_a0[4] ),
    .B1(\mul_wb.reg_a0[5] ),
    .C1(_3426_),
    .X(_3428_));
 sky130_fd_sc_hd__and2_2 _3858_ (.A(_3427_),
    .B(_3428_),
    .X(_3429_));
 sky130_fd_sc_hd__xor2_2 _3859_ (.A(\mul_wb.reg_a0[4] ),
    .B(_3426_),
    .X(_3430_));
 sky130_fd_sc_hd__xnor2_2 _3860_ (.A(\mul_wb.reg_a0[4] ),
    .B(_3426_),
    .Y(_3431_));
 sky130_fd_sc_hd__a21o_1 _3861_ (.A1(_3427_),
    .A2(_3428_),
    .B1(_3430_),
    .X(_3432_));
 sky130_fd_sc_hd__a211oi_2 _3862_ (.A1(_3427_),
    .A2(_3428_),
    .B1(_3430_),
    .C1(_3424_),
    .Y(_3433_));
 sky130_fd_sc_hd__and3_1 _3863_ (.A(net272),
    .B(_3421_),
    .C(_3433_),
    .X(_3434_));
 sky130_fd_sc_hd__and3_1 _3864_ (.A(_3412_),
    .B(_3419_),
    .C(_3434_),
    .X(_3435_));
 sky130_fd_sc_hd__nand2_1 _3865_ (.A(\mul_wb.lob_4.L[2] ),
    .B(_3388_),
    .Y(_3436_));
 sky130_fd_sc_hd__nand3_1 _3866_ (.A(\mul_wb.lob_4.L[3] ),
    .B(_3389_),
    .C(net250),
    .Y(_3437_));
 sky130_fd_sc_hd__a21oi_1 _3867_ (.A1(_3436_),
    .A2(_3437_),
    .B1(net248),
    .Y(_3438_));
 sky130_fd_sc_hd__a32o_1 _3868_ (.A1(\mul_wb.lob_4.L[7] ),
    .A2(_3407_),
    .A3(_3408_),
    .B1(\mul_wb.lob_4.L[5] ),
    .B2(net246),
    .X(_3439_));
 sky130_fd_sc_hd__a32o_1 _3869_ (.A1(_3384_),
    .A2(_3399_),
    .A3(_3439_),
    .B1(net248),
    .B2(\mul_wb.lob_4.L[1] ),
    .X(_3440_));
 sky130_fd_sc_hd__nor2_1 _3870_ (.A(_3388_),
    .B(net248),
    .Y(_3441_));
 sky130_fd_sc_hd__nand2_2 _3871_ (.A(_3389_),
    .B(_3396_),
    .Y(_3442_));
 sky130_fd_sc_hd__a21oi_2 _3872_ (.A1(_3381_),
    .A2(_3382_),
    .B1(net250),
    .Y(_3443_));
 sky130_fd_sc_hd__a2111oi_4 _3873_ (.A1(_3381_),
    .A2(_3382_),
    .B1(_3388_),
    .C1(net250),
    .D1(net248),
    .Y(_3444_));
 sky130_fd_sc_hd__a2111o_2 _3874_ (.A1(_3381_),
    .A2(_3382_),
    .B1(_3388_),
    .C1(net250),
    .D1(net248),
    .X(_3445_));
 sky130_fd_sc_hd__nor4_4 _3875_ (.A(net246),
    .B(_3405_),
    .C(_3408_),
    .D(_3415_),
    .Y(_3446_));
 sky130_fd_sc_hd__or4_1 _3876_ (.A(net246),
    .B(_3405_),
    .C(_3408_),
    .D(_3415_),
    .X(_3447_));
 sky130_fd_sc_hd__nor2_2 _3877_ (.A(_3417_),
    .B(_3429_),
    .Y(_3448_));
 sky130_fd_sc_hd__nand2_1 _3878_ (.A(net273),
    .B(_3424_),
    .Y(_3449_));
 sky130_fd_sc_hd__inv_2 _3879_ (.A(_3449_),
    .Y(_3450_));
 sky130_fd_sc_hd__and4_1 _3880_ (.A(_3431_),
    .B(_3446_),
    .C(_3448_),
    .D(_3450_),
    .X(_3451_));
 sky130_fd_sc_hd__and3_1 _3881_ (.A(\mul_wb.lob_4.L[6] ),
    .B(_3402_),
    .C(_3405_),
    .X(_3452_));
 sky130_fd_sc_hd__and4_1 _3882_ (.A(\mul_wb.lob_4.L[8] ),
    .B(_3407_),
    .C(_3409_),
    .D(_3415_),
    .X(_3453_));
 sky130_fd_sc_hd__o31a_1 _3883_ (.A1(_3451_),
    .A2(_3452_),
    .A3(_3453_),
    .B1(_3444_),
    .X(_3454_));
 sky130_fd_sc_hd__o41ai_4 _3884_ (.A1(_3435_),
    .A2(_3438_),
    .A3(_3440_),
    .A4(_3454_),
    .B1(\mul_wb.lob_4.A[0] ),
    .Y(_3455_));
 sky130_fd_sc_hd__a2111o_1 _3885_ (.A1(_3381_),
    .A2(_3382_),
    .B1(_3388_),
    .C1(net250),
    .D1(_3401_),
    .X(_3456_));
 sky130_fd_sc_hd__and3_1 _3886_ (.A(_3384_),
    .B(_3399_),
    .C(_3402_),
    .X(_3457_));
 sky130_fd_sc_hd__nor3_1 _3887_ (.A(_3408_),
    .B(_3415_),
    .C(_3418_),
    .Y(_3458_));
 sky130_fd_sc_hd__nand2_1 _3888_ (.A(\mul_wb.lob_4.A[0] ),
    .B(net266),
    .Y(_3459_));
 sky130_fd_sc_hd__xor2_2 _3889_ (.A(\mul_wb.reg_a0[1] ),
    .B(_3459_),
    .X(_3460_));
 sky130_fd_sc_hd__and4_1 _3890_ (.A(\mul_wb.lob_4.A[0] ),
    .B(net274),
    .C(_3416_),
    .D(_3430_),
    .X(_3461_));
 sky130_fd_sc_hd__and3b_1 _3891_ (.A_N(net250),
    .B(\mul_wb.lob_4.L[4] ),
    .C(\mul_wb.lob_4.A[0] ),
    .X(_3462_));
 sky130_fd_sc_hd__and3_1 _3892_ (.A(_3383_),
    .B(_3441_),
    .C(_3462_),
    .X(_3463_));
 sky130_fd_sc_hd__or4_1 _3893_ (.A(_3363_),
    .B(_3365_),
    .C(_3421_),
    .D(_3460_),
    .X(_3464_));
 sky130_fd_sc_hd__or4b_1 _3894_ (.A(_3363_),
    .B(_3421_),
    .C(_3424_),
    .D_N(_3460_),
    .X(_3465_));
 sky130_fd_sc_hd__or4_1 _3895_ (.A(_3415_),
    .B(_3417_),
    .C(_3432_),
    .D(_3465_),
    .X(_3466_));
 sky130_fd_sc_hd__or4_2 _3896_ (.A(_3364_),
    .B(_3400_),
    .C(_3411_),
    .D(_3466_),
    .X(_3467_));
 sky130_fd_sc_hd__and4_1 _3897_ (.A(\mul_wb.lob_4.A[0] ),
    .B(net275),
    .C(_3418_),
    .D(_3429_),
    .X(_3468_));
 sky130_fd_sc_hd__and3_1 _3898_ (.A(_3444_),
    .B(_3446_),
    .C(_3468_),
    .X(_3469_));
 sky130_fd_sc_hd__and4_1 _3899_ (.A(\mul_wb.lob_4.A[0] ),
    .B(\mul_wb.lob_4.L[9] ),
    .C(_3406_),
    .D(_3458_),
    .X(_3470_));
 sky130_fd_sc_hd__a211o_1 _3900_ (.A1(_3457_),
    .A2(_3470_),
    .B1(_3469_),
    .C1(_3463_),
    .X(_3471_));
 sky130_fd_sc_hd__nand2_1 _3901_ (.A(_3418_),
    .B(_3433_),
    .Y(_3472_));
 sky130_fd_sc_hd__nor4_1 _3902_ (.A(_3445_),
    .B(_3447_),
    .C(_3464_),
    .D(_3472_),
    .Y(_3473_));
 sky130_fd_sc_hd__a311oi_4 _3903_ (.A1(_3412_),
    .A2(_3448_),
    .A3(_3461_),
    .B1(_3471_),
    .C1(net228),
    .Y(_3474_));
 sky130_fd_sc_hd__and3_4 _3904_ (.A(_3455_),
    .B(_3467_),
    .C(_3474_),
    .X(_3475_));
 sky130_fd_sc_hd__or4_4 _3905_ (.A(\mul_wb.reg_b0[1] ),
    .B(\mul_wb.lob_4.B[0] ),
    .C(\mul_wb.reg_b0[2] ),
    .D(\mul_wb.reg_b0[3] ),
    .X(_3476_));
 sky130_fd_sc_hd__or4_4 _3906_ (.A(\mul_wb.reg_b0[4] ),
    .B(\mul_wb.reg_b0[5] ),
    .C(\mul_wb.reg_b0[6] ),
    .D(\mul_wb.reg_b0[7] ),
    .X(_3477_));
 sky130_fd_sc_hd__or2_1 _3907_ (.A(\mul_wb.reg_b0[8] ),
    .B(\mul_wb.reg_b0[9] ),
    .X(_3478_));
 sky130_fd_sc_hd__or4_2 _3908_ (.A(\mul_wb.reg_b0[8] ),
    .B(\mul_wb.reg_b0[9] ),
    .C(\mul_wb.reg_b0[10] ),
    .D(\mul_wb.reg_b0[11] ),
    .X(_3479_));
 sky130_fd_sc_hd__or2_1 _3909_ (.A(\mul_wb.reg_b0[12] ),
    .B(\mul_wb.reg_b0[13] ),
    .X(_3480_));
 sky130_fd_sc_hd__or4_1 _3910_ (.A(_3476_),
    .B(_3477_),
    .C(_3479_),
    .D(_3480_),
    .X(_3481_));
 sky130_fd_sc_hd__o41a_2 _3911_ (.A1(_3476_),
    .A2(_3477_),
    .A3(_3479_),
    .A4(_3480_),
    .B1(net267),
    .X(_3482_));
 sky130_fd_sc_hd__xor2_4 _3912_ (.A(\mul_wb.reg_b0[14] ),
    .B(_3482_),
    .X(_3483_));
 sky130_fd_sc_hd__xnor2_2 _3913_ (.A(\mul_wb.reg_b0[14] ),
    .B(_3482_),
    .Y(_3484_));
 sky130_fd_sc_hd__o31a_2 _3914_ (.A1(_3476_),
    .A2(_3477_),
    .A3(_3478_),
    .B1(\mul_wb.reg_b0[15] ),
    .X(_3485_));
 sky130_fd_sc_hd__o41a_2 _3915_ (.A1(\mul_wb.reg_b0[10] ),
    .A2(_3476_),
    .A3(_3477_),
    .A4(_3478_),
    .B1(net267),
    .X(_3486_));
 sky130_fd_sc_hd__xor2_4 _3916_ (.A(\mul_wb.reg_b0[11] ),
    .B(_3486_),
    .X(_3487_));
 sky130_fd_sc_hd__xor2_4 _3917_ (.A(\mul_wb.reg_b0[10] ),
    .B(_3485_),
    .X(_3488_));
 sky130_fd_sc_hd__xnor2_2 _3918_ (.A(\mul_wb.reg_b0[10] ),
    .B(_3485_),
    .Y(_3489_));
 sky130_fd_sc_hd__or3b_1 _3919_ (.A(_3487_),
    .B(_3489_),
    .C_N(\mul_wb.lob_4.L[5] ),
    .X(_3490_));
 sky130_fd_sc_hd__nand2_1 _3920_ (.A(\mul_wb.lob_4.L[4] ),
    .B(_3487_),
    .Y(_3491_));
 sky130_fd_sc_hd__o31a_1 _3921_ (.A1(_3476_),
    .A2(_3477_),
    .A3(_3479_),
    .B1(net267),
    .X(_3492_));
 sky130_fd_sc_hd__xor2_2 _3922_ (.A(\mul_wb.reg_b0[12] ),
    .B(_3492_),
    .X(_3493_));
 sky130_fd_sc_hd__o41a_4 _3923_ (.A1(\mul_wb.reg_b0[12] ),
    .A2(_3476_),
    .A3(_3477_),
    .A4(_3479_),
    .B1(net267),
    .X(_3494_));
 sky130_fd_sc_hd__xor2_4 _3924_ (.A(\mul_wb.reg_b0[13] ),
    .B(_3494_),
    .X(_3495_));
 sky130_fd_sc_hd__xnor2_4 _3925_ (.A(\mul_wb.reg_b0[13] ),
    .B(_3494_),
    .Y(_3496_));
 sky130_fd_sc_hd__nor2_1 _3926_ (.A(net243),
    .B(_3495_),
    .Y(_3497_));
 sky130_fd_sc_hd__nor3b_4 _3927_ (.A(net969),
    .B(_3481_),
    .C_N(net267),
    .Y(_3498_));
 sky130_fd_sc_hd__and2_1 _3928_ (.A(net243),
    .B(_3496_),
    .X(_3499_));
 sky130_fd_sc_hd__a21oi_1 _3929_ (.A1(_3490_),
    .A2(_3491_),
    .B1(net243),
    .Y(_3500_));
 sky130_fd_sc_hd__a211o_1 _3930_ (.A1(\mul_wb.lob_4.L[3] ),
    .A2(net243),
    .B1(_3495_),
    .C1(_3500_),
    .X(_3501_));
 sky130_fd_sc_hd__nor2_1 _3931_ (.A(_3487_),
    .B(net243),
    .Y(_3502_));
 sky130_fd_sc_hd__nor4_4 _3932_ (.A(_3487_),
    .B(_3488_),
    .C(net243),
    .D(_3495_),
    .Y(_3503_));
 sky130_fd_sc_hd__o21ai_2 _3933_ (.A1(_3476_),
    .A2(_3477_),
    .B1(net267),
    .Y(_3504_));
 sky130_fd_sc_hd__o31a_2 _3934_ (.A1(\mul_wb.reg_b0[8] ),
    .A2(_3476_),
    .A3(_3477_),
    .B1(net267),
    .X(_3505_));
 sky130_fd_sc_hd__xor2_4 _3935_ (.A(\mul_wb.reg_b0[9] ),
    .B(_3505_),
    .X(_3506_));
 sky130_fd_sc_hd__xnor2_4 _3936_ (.A(\mul_wb.reg_b0[8] ),
    .B(_3504_),
    .Y(_3507_));
 sky130_fd_sc_hd__nor2_1 _3937_ (.A(_3506_),
    .B(_3507_),
    .Y(_3508_));
 sky130_fd_sc_hd__o31a_2 _3938_ (.A1(\mul_wb.reg_b0[4] ),
    .A2(\mul_wb.reg_b0[5] ),
    .A3(_3476_),
    .B1(net267),
    .X(_3509_));
 sky130_fd_sc_hd__o41a_2 _3939_ (.A1(\mul_wb.reg_b0[4] ),
    .A2(\mul_wb.reg_b0[5] ),
    .A3(\mul_wb.reg_b0[6] ),
    .A4(_3476_),
    .B1(net267),
    .X(_3510_));
 sky130_fd_sc_hd__xor2_4 _3940_ (.A(\mul_wb.reg_b0[7] ),
    .B(_3510_),
    .X(_3511_));
 sky130_fd_sc_hd__and4_1 _3941_ (.A(\mul_wb.lob_4.L[8] ),
    .B(net244),
    .C(_3503_),
    .D(_3511_),
    .X(_3512_));
 sky130_fd_sc_hd__nor2_4 _3942_ (.A(_3483_),
    .B(_3498_),
    .Y(_3513_));
 sky130_fd_sc_hd__and2_1 _3943_ (.A(_3503_),
    .B(_3513_),
    .X(_3514_));
 sky130_fd_sc_hd__xor2_4 _3944_ (.A(\mul_wb.reg_b0[6] ),
    .B(_3509_),
    .X(_3515_));
 sky130_fd_sc_hd__inv_2 _3945_ (.A(_3515_),
    .Y(_3516_));
 sky130_fd_sc_hd__and3b_1 _3946_ (.A_N(_3511_),
    .B(_3515_),
    .C(\mul_wb.lob_4.L[9] ),
    .X(_3517_));
 sky130_fd_sc_hd__and3_1 _3947_ (.A(_3503_),
    .B(_3513_),
    .C(_3517_),
    .X(_3518_));
 sky130_fd_sc_hd__o21a_1 _3948_ (.A1(_3512_),
    .A2(_3518_),
    .B1(_3508_),
    .X(_3519_));
 sky130_fd_sc_hd__o31a_2 _3949_ (.A1(\mul_wb.reg_b0[1] ),
    .A2(\mul_wb.lob_4.B[0] ),
    .A3(\mul_wb.reg_b0[2] ),
    .B1(net267),
    .X(_3520_));
 sky130_fd_sc_hd__xor2_4 _3950_ (.A(\mul_wb.reg_b0[3] ),
    .B(_3520_),
    .X(_3521_));
 sky130_fd_sc_hd__o21ai_2 _3951_ (.A1(\mul_wb.reg_b0[4] ),
    .A2(_3476_),
    .B1(net267),
    .Y(_3522_));
 sky130_fd_sc_hd__xnor2_4 _3952_ (.A(\mul_wb.reg_b0[5] ),
    .B(_3522_),
    .Y(_3523_));
 sky130_fd_sc_hd__a21oi_1 _3953_ (.A1(net267),
    .A2(_3476_),
    .B1(\mul_wb.reg_b0[4] ),
    .Y(_3524_));
 sky130_fd_sc_hd__and3_1 _3954_ (.A(net267),
    .B(\mul_wb.reg_b0[4] ),
    .C(_3476_),
    .X(_3525_));
 sky130_fd_sc_hd__nor2_4 _3955_ (.A(_3524_),
    .B(_3525_),
    .Y(_3526_));
 sky130_fd_sc_hd__inv_2 _3956_ (.A(_3526_),
    .Y(_3527_));
 sky130_fd_sc_hd__nor2_1 _3957_ (.A(_3523_),
    .B(_3526_),
    .Y(_3528_));
 sky130_fd_sc_hd__nor2_1 _3958_ (.A(_3507_),
    .B(_3511_),
    .Y(_3529_));
 sky130_fd_sc_hd__nor4_1 _3959_ (.A(_3506_),
    .B(_3507_),
    .C(_3511_),
    .D(_3515_),
    .Y(_3530_));
 sky130_fd_sc_hd__and2_1 _3960_ (.A(_3528_),
    .B(net240),
    .X(_3531_));
 sky130_fd_sc_hd__o21ai_2 _3961_ (.A1(\mul_wb.reg_b0[1] ),
    .A2(\mul_wb.lob_4.B[0] ),
    .B1(net267),
    .Y(_3532_));
 sky130_fd_sc_hd__xnor2_4 _3962_ (.A(\mul_wb.reg_b0[2] ),
    .B(_3532_),
    .Y(_3533_));
 sky130_fd_sc_hd__nand2_2 _3963_ (.A(\mul_wb.lob_4.B[0] ),
    .B(net267),
    .Y(_3534_));
 sky130_fd_sc_hd__xnor2_4 _3964_ (.A(\mul_wb.reg_b0[1] ),
    .B(_3534_),
    .Y(_3535_));
 sky130_fd_sc_hd__nor2_1 _3965_ (.A(_3533_),
    .B(_3535_),
    .Y(_3536_));
 sky130_fd_sc_hd__a22o_1 _3966_ (.A1(\mul_wb.lob_4.L[13] ),
    .A2(_3533_),
    .B1(_3536_),
    .B2(net268),
    .X(_3537_));
 sky130_fd_sc_hd__and4b_1 _3967_ (.A_N(_3521_),
    .B(_3528_),
    .C(_3530_),
    .D(_3537_),
    .X(_3538_));
 sky130_fd_sc_hd__and3b_1 _3968_ (.A_N(_3506_),
    .B(_3507_),
    .C(\mul_wb.lob_4.L[7] ),
    .X(_3539_));
 sky130_fd_sc_hd__o21a_1 _3969_ (.A1(_3538_),
    .A2(_3539_),
    .B1(_3514_),
    .X(_3540_));
 sky130_fd_sc_hd__nand2_1 _3970_ (.A(net244),
    .B(_3496_),
    .Y(_3541_));
 sky130_fd_sc_hd__inv_2 _3971_ (.A(_3541_),
    .Y(_3542_));
 sky130_fd_sc_hd__nor4_2 _3972_ (.A(_3483_),
    .B(_3487_),
    .C(net243),
    .D(_3495_),
    .Y(_3543_));
 sky130_fd_sc_hd__nor2_1 _3973_ (.A(_3488_),
    .B(_3506_),
    .Y(_3544_));
 sky130_fd_sc_hd__nor4_1 _3974_ (.A(_3488_),
    .B(_3506_),
    .C(_3507_),
    .D(_3511_),
    .Y(_3545_));
 sky130_fd_sc_hd__and2_1 _3975_ (.A(net239),
    .B(_3545_),
    .X(_3546_));
 sky130_fd_sc_hd__a32o_1 _3976_ (.A1(net273),
    .A2(_3521_),
    .A3(_3528_),
    .B1(_3523_),
    .B2(net275),
    .X(_3547_));
 sky130_fd_sc_hd__and2_1 _3977_ (.A(\mul_wb.lob_4.L[1] ),
    .B(_3483_),
    .X(_3548_));
 sky130_fd_sc_hd__a41o_1 _3978_ (.A1(\mul_wb.lob_4.L[6] ),
    .A2(net244),
    .A3(_3503_),
    .A4(_3506_),
    .B1(_3548_),
    .X(_3549_));
 sky130_fd_sc_hd__a31o_1 _3979_ (.A1(_3516_),
    .A2(_3546_),
    .A3(_3547_),
    .B1(_3549_),
    .X(_3550_));
 sky130_fd_sc_hd__o21a_1 _3980_ (.A1(\mul_wb.lob_4.L[2] ),
    .A2(_3496_),
    .B1(net244),
    .X(_3551_));
 sky130_fd_sc_hd__a2111o_1 _3981_ (.A1(_3501_),
    .A2(_3551_),
    .B1(_3550_),
    .C1(_3540_),
    .D1(_3519_),
    .X(_3552_));
 sky130_fd_sc_hd__nor4_2 _3982_ (.A(_3483_),
    .B(_3498_),
    .C(_3506_),
    .D(_3507_),
    .Y(_3553_));
 sky130_fd_sc_hd__nor2_1 _3983_ (.A(_3515_),
    .B(_3523_),
    .Y(_3554_));
 sky130_fd_sc_hd__and4b_1 _3984_ (.A_N(_3511_),
    .B(_3526_),
    .C(net274),
    .D(\mul_wb.lob_4.B[0] ),
    .X(_3555_));
 sky130_fd_sc_hd__nor4_1 _3985_ (.A(_3515_),
    .B(_3521_),
    .C(_3523_),
    .D(_3526_),
    .Y(_3556_));
 sky130_fd_sc_hd__and2_1 _3986_ (.A(_3529_),
    .B(_3556_),
    .X(_3557_));
 sky130_fd_sc_hd__and3_1 _3987_ (.A(_3535_),
    .B(net239),
    .C(_3544_),
    .X(_3558_));
 sky130_fd_sc_hd__and3b_1 _3988_ (.A_N(_3533_),
    .B(\mul_wb.lob_4.B[0] ),
    .C(net270),
    .X(_3559_));
 sky130_fd_sc_hd__and4_1 _3989_ (.A(_3503_),
    .B(_3553_),
    .C(_3554_),
    .D(_3555_),
    .X(_3560_));
 sky130_fd_sc_hd__a31o_1 _3990_ (.A1(_3557_),
    .A2(_3558_),
    .A3(_3559_),
    .B1(_3560_),
    .X(_3561_));
 sky130_fd_sc_hd__a21oi_1 _3991_ (.A1(net705),
    .A2(_3552_),
    .B1(_3561_),
    .Y(_3562_));
 sky130_fd_sc_hd__nor2_1 _3992_ (.A(net177),
    .B(net176),
    .Y(\mul_wb.P_[0] ));
 sky130_fd_sc_hd__and4bb_1 _3993_ (.A_N(_3415_),
    .B_N(_3432_),
    .C(_3418_),
    .D(_3424_),
    .X(_3563_));
 sky130_fd_sc_hd__or4b_1 _3994_ (.A(_3366_),
    .B(_3400_),
    .C(_3411_),
    .D_N(_3563_),
    .X(_3564_));
 sky130_fd_sc_hd__and3_1 _3995_ (.A(_3417_),
    .B(net241),
    .C(_3446_),
    .X(_3565_));
 sky130_fd_sc_hd__and4_1 _3996_ (.A(net275),
    .B(_3417_),
    .C(net241),
    .D(_3446_),
    .X(_3566_));
 sky130_fd_sc_hd__nor2_1 _3997_ (.A(_3384_),
    .B(_3400_),
    .Y(_3567_));
 sky130_fd_sc_hd__and3_1 _3998_ (.A(_3389_),
    .B(_3390_),
    .C(_3396_),
    .X(_3568_));
 sky130_fd_sc_hd__nand2_1 _3999_ (.A(\mul_wb.lob_4.L[4] ),
    .B(_3568_),
    .Y(_3569_));
 sky130_fd_sc_hd__nor2_2 _4000_ (.A(_3389_),
    .B(net248),
    .Y(_3570_));
 sky130_fd_sc_hd__a22oi_1 _4001_ (.A1(\mul_wb.lob_4.L[2] ),
    .A2(net249),
    .B1(_3570_),
    .B2(\mul_wb.lob_4.L[3] ),
    .Y(_3571_));
 sky130_fd_sc_hd__nand3_1 _4002_ (.A(_3443_),
    .B(_3446_),
    .C(_3448_),
    .Y(_3572_));
 sky130_fd_sc_hd__and3_1 _4003_ (.A(_3389_),
    .B(_3396_),
    .C(_3430_),
    .X(_3573_));
 sky130_fd_sc_hd__nand2_1 _4004_ (.A(net273),
    .B(_3573_),
    .Y(_3574_));
 sky130_fd_sc_hd__nand3_1 _4005_ (.A(\mul_wb.lob_4.L[6] ),
    .B(net246),
    .C(net241),
    .Y(_3575_));
 sky130_fd_sc_hd__or3_1 _4006_ (.A(net248),
    .B(_3397_),
    .C(_3406_),
    .X(_3576_));
 sky130_fd_sc_hd__nor2_2 _4007_ (.A(_3456_),
    .B(_3576_),
    .Y(_3577_));
 sky130_fd_sc_hd__and3_1 _4008_ (.A(_3399_),
    .B(_3410_),
    .C(_3415_),
    .X(_3578_));
 sky130_fd_sc_hd__a32o_1 _4009_ (.A1(net268),
    .A2(_3422_),
    .A3(_3433_),
    .B1(_3429_),
    .B2(net274),
    .X(_3579_));
 sky130_fd_sc_hd__or4_1 _4010_ (.A(_3422_),
    .B(_3445_),
    .C(_3447_),
    .D(_3472_),
    .X(_3580_));
 sky130_fd_sc_hd__nand4_1 _4011_ (.A(\mul_wb.lob_4.L[8] ),
    .B(_3407_),
    .C(_3408_),
    .D(net241),
    .Y(_3581_));
 sky130_fd_sc_hd__a32oi_1 _4012_ (.A1(_3412_),
    .A2(_3419_),
    .A3(_3579_),
    .B1(_3567_),
    .B2(\mul_wb.lob_4.L[5] ),
    .Y(_3582_));
 sky130_fd_sc_hd__a31o_1 _4013_ (.A1(_3569_),
    .A2(_3581_),
    .A3(_3582_),
    .B1(_3460_),
    .X(_3583_));
 sky130_fd_sc_hd__o221a_1 _4014_ (.A1(_3572_),
    .A2(_3574_),
    .B1(_3580_),
    .B2(_3365_),
    .C1(_3564_),
    .X(_3584_));
 sky130_fd_sc_hd__a221oi_1 _4015_ (.A1(\mul_wb.lob_4.L[7] ),
    .A2(_3577_),
    .B1(_3578_),
    .B2(\mul_wb.lob_4.L[9] ),
    .C1(_3566_),
    .Y(_3585_));
 sky130_fd_sc_hd__a41o_1 _4016_ (.A1(_3571_),
    .A2(_3575_),
    .A3(_3584_),
    .A4(_3585_),
    .B1(_3460_),
    .X(_3586_));
 sky130_fd_sc_hd__and2_2 _4017_ (.A(_3583_),
    .B(_3586_),
    .X(_3587_));
 sky130_fd_sc_hd__and3_1 _4018_ (.A(_3521_),
    .B(_3528_),
    .C(net240),
    .X(_3588_));
 sky130_fd_sc_hd__nor2_2 _4019_ (.A(net245),
    .B(_3496_),
    .Y(_3589_));
 sky130_fd_sc_hd__and3_1 _4020_ (.A(_3515_),
    .B(_3543_),
    .C(net238),
    .X(_3590_));
 sky130_fd_sc_hd__and4_1 _4021_ (.A(net275),
    .B(_3515_),
    .C(net239),
    .D(_3545_),
    .X(_3591_));
 sky130_fd_sc_hd__and3_2 _4022_ (.A(_3503_),
    .B(_3506_),
    .C(_3513_),
    .X(_3592_));
 sky130_fd_sc_hd__and3_1 _4023_ (.A(_3503_),
    .B(_3511_),
    .C(_3553_),
    .X(_3593_));
 sky130_fd_sc_hd__and3_1 _4024_ (.A(net269),
    .B(_3503_),
    .C(_3513_),
    .X(_3594_));
 sky130_fd_sc_hd__and4bb_1 _4025_ (.A_N(_3521_),
    .B_N(_3533_),
    .C(_3594_),
    .D(_3531_),
    .X(_3595_));
 sky130_fd_sc_hd__nor4_1 _4026_ (.A(_3487_),
    .B(net243),
    .C(_3515_),
    .D(_3523_),
    .Y(_3596_));
 sky130_fd_sc_hd__and3_1 _4027_ (.A(net244),
    .B(_3496_),
    .C(_3526_),
    .X(_3597_));
 sky130_fd_sc_hd__a32o_1 _4028_ (.A1(net271),
    .A2(_3533_),
    .A3(_3557_),
    .B1(\mul_wb.lob_4.L[8] ),
    .B2(_3507_),
    .X(_3598_));
 sky130_fd_sc_hd__and4_1 _4029_ (.A(_3503_),
    .B(_3513_),
    .C(_3523_),
    .D(net240),
    .X(_3599_));
 sky130_fd_sc_hd__and3_2 _4030_ (.A(_3487_),
    .B(_3497_),
    .C(_3513_),
    .X(_3600_));
 sky130_fd_sc_hd__and3_1 _4031_ (.A(net244),
    .B(net243),
    .C(_3496_),
    .X(_3601_));
 sky130_fd_sc_hd__and3_1 _4032_ (.A(\mul_wb.lob_4.L[4] ),
    .B(_3535_),
    .C(_3601_),
    .X(_3602_));
 sky130_fd_sc_hd__and3_1 _4033_ (.A(\mul_wb.lob_4.L[9] ),
    .B(_3511_),
    .C(_3535_),
    .X(_3603_));
 sky130_fd_sc_hd__and3_1 _4034_ (.A(_3503_),
    .B(_3553_),
    .C(_3603_),
    .X(_3604_));
 sky130_fd_sc_hd__a311o_1 _4035_ (.A1(\mul_wb.lob_4.L[5] ),
    .A2(_3535_),
    .A3(_3600_),
    .B1(_3602_),
    .C1(_3604_),
    .X(_3605_));
 sky130_fd_sc_hd__and2_1 _4036_ (.A(_3503_),
    .B(net240),
    .X(_3606_));
 sky130_fd_sc_hd__a41o_1 _4037_ (.A1(net274),
    .A2(_3513_),
    .A3(_3523_),
    .A4(_3606_),
    .B1(_3591_),
    .X(_3607_));
 sky130_fd_sc_hd__a221oi_4 _4038_ (.A1(_3558_),
    .A2(_3598_),
    .B1(_3607_),
    .B2(_3535_),
    .C1(_3605_),
    .Y(_3608_));
 sky130_fd_sc_hd__a32o_1 _4039_ (.A1(\mul_wb.lob_4.L[6] ),
    .A2(_3488_),
    .A3(net239),
    .B1(\mul_wb.lob_4.L[2] ),
    .B2(net245),
    .X(_3609_));
 sky130_fd_sc_hd__a221o_1 _4040_ (.A1(\mul_wb.lob_4.L[3] ),
    .A2(_3589_),
    .B1(_3592_),
    .B2(\mul_wb.lob_4.L[7] ),
    .C1(_3609_),
    .X(_3610_));
 sky130_fd_sc_hd__and4_1 _4041_ (.A(net273),
    .B(net238),
    .C(_3596_),
    .D(_3597_),
    .X(_3611_));
 sky130_fd_sc_hd__a41o_1 _4042_ (.A1(net272),
    .A2(_3514_),
    .A3(_3521_),
    .A4(_3531_),
    .B1(_3611_),
    .X(_3612_));
 sky130_fd_sc_hd__o31ai_4 _4043_ (.A1(_3595_),
    .A2(_3610_),
    .A3(_3612_),
    .B1(_3535_),
    .Y(_3613_));
 sky130_fd_sc_hd__and2_4 _4044_ (.A(_3608_),
    .B(_3613_),
    .X(_3614_));
 sky130_fd_sc_hd__o22ai_1 _4045_ (.A1(net176),
    .A2(net174),
    .B1(_3614_),
    .B2(net177),
    .Y(_3615_));
 sky130_fd_sc_hd__or4_1 _4046_ (.A(net177),
    .B(net176),
    .C(net174),
    .D(_3614_),
    .X(_3616_));
 sky130_fd_sc_hd__inv_2 _4047_ (.A(_3616_),
    .Y(_3617_));
 sky130_fd_sc_hd__nand2_1 _4048_ (.A(_3615_),
    .B(_3616_),
    .Y(_3618_));
 sky130_fd_sc_hd__xor2_1 _4049_ (.A(\mul_wb.reg_a0[15] ),
    .B(net697),
    .X(_3619_));
 sky130_fd_sc_hd__xnor2_4 _4050_ (.A(net703),
    .B(net267),
    .Y(_3620_));
 sky130_fd_sc_hd__nand2_1 _4051_ (.A(\mul_wb.P_[0] ),
    .B(net252),
    .Y(_3621_));
 sky130_fd_sc_hd__xor2_1 _4052_ (.A(_3618_),
    .B(_3621_),
    .X(\mul_wb.reg_p[1] ));
 sky130_fd_sc_hd__or2_1 _4053_ (.A(\mul_wb.P_[0] ),
    .B(_3615_),
    .X(_3622_));
 sky130_fd_sc_hd__nand2_1 _4054_ (.A(net252),
    .B(_3622_),
    .Y(_3623_));
 sky130_fd_sc_hd__or2_1 _4055_ (.A(net174),
    .B(_3614_),
    .X(_3624_));
 sky130_fd_sc_hd__nor2_1 _4056_ (.A(\mul_wb.P_[0] ),
    .B(_3624_),
    .Y(_3625_));
 sky130_fd_sc_hd__and3_1 _4057_ (.A(_3507_),
    .B(net239),
    .C(_3544_),
    .X(_3626_));
 sky130_fd_sc_hd__a22o_1 _4058_ (.A1(net274),
    .A2(_3590_),
    .B1(_3626_),
    .B2(\mul_wb.lob_4.L[9] ),
    .X(_3627_));
 sky130_fd_sc_hd__a32o_1 _4059_ (.A1(net271),
    .A2(_3514_),
    .A3(_3588_),
    .B1(_3592_),
    .B2(\mul_wb.lob_4.L[8] ),
    .X(_3628_));
 sky130_fd_sc_hd__nand2_1 _4060_ (.A(\mul_wb.lob_4.L[5] ),
    .B(net243),
    .Y(_3629_));
 sky130_fd_sc_hd__or4b_1 _4061_ (.A(_3487_),
    .B(_3489_),
    .C(net243),
    .D_N(\mul_wb.lob_4.L[7] ),
    .X(_3630_));
 sky130_fd_sc_hd__a21oi_1 _4062_ (.A1(_3629_),
    .A2(_3630_),
    .B1(_3495_),
    .Y(_3631_));
 sky130_fd_sc_hd__and3b_1 _4063_ (.A_N(net243),
    .B(_3496_),
    .C(_3487_),
    .X(_3632_));
 sky130_fd_sc_hd__a22o_1 _4064_ (.A1(\mul_wb.lob_4.L[4] ),
    .A2(_3495_),
    .B1(_3632_),
    .B2(\mul_wb.lob_4.L[6] ),
    .X(_3633_));
 sky130_fd_sc_hd__o21a_1 _4065_ (.A1(_3631_),
    .A2(_3633_),
    .B1(net244),
    .X(_3634_));
 sky130_fd_sc_hd__and4_1 _4066_ (.A(net272),
    .B(net238),
    .C(_3596_),
    .D(_3597_),
    .X(_3635_));
 sky130_fd_sc_hd__and3b_1 _4067_ (.A_N(_3506_),
    .B(net269),
    .C(_3489_),
    .X(_3636_));
 sky130_fd_sc_hd__and2_1 _4068_ (.A(\mul_wb.lob_4.L[3] ),
    .B(_3483_),
    .X(_3637_));
 sky130_fd_sc_hd__a41o_1 _4069_ (.A1(_3529_),
    .A2(net239),
    .A3(_3556_),
    .A4(_3636_),
    .B1(_3637_),
    .X(_3638_));
 sky130_fd_sc_hd__and4_1 _4070_ (.A(net275),
    .B(_3503_),
    .C(_3511_),
    .D(_3553_),
    .X(_3639_));
 sky130_fd_sc_hd__a2111o_1 _4071_ (.A1(net273),
    .A2(_3599_),
    .B1(_3635_),
    .C1(_3638_),
    .D1(_3639_),
    .X(_3640_));
 sky130_fd_sc_hd__o41ai_2 _4072_ (.A1(_3627_),
    .A2(_3628_),
    .A3(_3634_),
    .A4(_3640_),
    .B1(_3533_),
    .Y(_3641_));
 sky130_fd_sc_hd__and3_1 _4073_ (.A(\mul_wb.lob_4.L[6] ),
    .B(_3383_),
    .C(_3399_),
    .X(_3642_));
 sky130_fd_sc_hd__a22o_1 _4074_ (.A1(\mul_wb.lob_4.L[9] ),
    .A2(_3408_),
    .B1(_3458_),
    .B2(net274),
    .X(_3643_));
 sky130_fd_sc_hd__and2_1 _4075_ (.A(\mul_wb.lob_4.L[8] ),
    .B(_3577_),
    .X(_3644_));
 sky130_fd_sc_hd__a32o_1 _4076_ (.A1(\mul_wb.lob_4.L[7] ),
    .A2(net246),
    .A3(_3443_),
    .B1(\mul_wb.lob_4.L[5] ),
    .B2(net250),
    .X(_3645_));
 sky130_fd_sc_hd__a32o_1 _4077_ (.A1(_3407_),
    .A2(net241),
    .A3(_3643_),
    .B1(_3578_),
    .B2(net275),
    .X(_3646_));
 sky130_fd_sc_hd__a221o_1 _4078_ (.A1(\mul_wb.lob_4.L[3] ),
    .A2(net249),
    .B1(_3441_),
    .B2(_3645_),
    .C1(_3642_),
    .X(_3647_));
 sky130_fd_sc_hd__o31ai_4 _4079_ (.A1(_3644_),
    .A2(_3646_),
    .A3(_3647_),
    .B1(_3421_),
    .Y(_3648_));
 sky130_fd_sc_hd__and4_1 _4080_ (.A(_3399_),
    .B(_3410_),
    .C(_3419_),
    .D(_3429_),
    .X(_3649_));
 sky130_fd_sc_hd__and3_1 _4081_ (.A(net273),
    .B(_3421_),
    .C(_3649_),
    .X(_3650_));
 sky130_fd_sc_hd__and4_1 _4082_ (.A(net270),
    .B(_3412_),
    .C(_3421_),
    .D(_3563_),
    .X(_3651_));
 sky130_fd_sc_hd__and3_1 _4083_ (.A(\mul_wb.lob_4.L[4] ),
    .B(_3421_),
    .C(_3570_),
    .X(_3652_));
 sky130_fd_sc_hd__or3b_1 _4084_ (.A(_3366_),
    .B(_3422_),
    .C_N(_3573_),
    .X(_3653_));
 sky130_fd_sc_hd__o21ba_1 _4085_ (.A1(_3572_),
    .A2(_3653_),
    .B1_N(_3652_),
    .X(_3654_));
 sky130_fd_sc_hd__or2_1 _4086_ (.A(_3364_),
    .B(_3580_),
    .X(_3655_));
 sky130_fd_sc_hd__and4bb_2 _4087_ (.A_N(_3650_),
    .B_N(_3651_),
    .C(_3654_),
    .D(_3655_),
    .X(_3656_));
 sky130_fd_sc_hd__and2_2 _4088_ (.A(_3648_),
    .B(_3656_),
    .X(_3657_));
 sky130_fd_sc_hd__or2_1 _4089_ (.A(net176),
    .B(net173),
    .X(_3658_));
 sky130_fd_sc_hd__nor3_1 _4090_ (.A(net177),
    .B(net210),
    .C(_3658_),
    .Y(_3659_));
 sky130_fd_sc_hd__o21a_1 _4091_ (.A1(net177),
    .A2(net210),
    .B1(_3658_),
    .X(_3660_));
 sky130_fd_sc_hd__or2_2 _4092_ (.A(_3659_),
    .B(_3660_),
    .X(_3661_));
 sky130_fd_sc_hd__nor2_1 _4093_ (.A(_3624_),
    .B(_3661_),
    .Y(_3662_));
 sky130_fd_sc_hd__xnor2_1 _4094_ (.A(_3625_),
    .B(_3661_),
    .Y(_3663_));
 sky130_fd_sc_hd__xnor2_1 _4095_ (.A(_3623_),
    .B(_3663_),
    .Y(\mul_wb.reg_p[2] ));
 sky130_fd_sc_hd__or2_1 _4096_ (.A(_3622_),
    .B(_3663_),
    .X(_3664_));
 sky130_fd_sc_hd__nand2_1 _4097_ (.A(net252),
    .B(_3664_),
    .Y(_3665_));
 sky130_fd_sc_hd__nor2_1 _4098_ (.A(net174),
    .B(net210),
    .Y(_3666_));
 sky130_fd_sc_hd__and2_1 _4099_ (.A(\mul_wb.lob_4.L[6] ),
    .B(net250),
    .X(_3667_));
 sky130_fd_sc_hd__nand2_1 _4100_ (.A(net270),
    .B(_3430_),
    .Y(_3668_));
 sky130_fd_sc_hd__inv_2 _4101_ (.A(_3668_),
    .Y(_3669_));
 sky130_fd_sc_hd__a41o_1 _4102_ (.A1(_3443_),
    .A2(_3446_),
    .A3(_3448_),
    .A4(_3669_),
    .B1(_3667_),
    .X(_3670_));
 sky130_fd_sc_hd__nor2_1 _4103_ (.A(_3425_),
    .B(_3442_),
    .Y(_3671_));
 sky130_fd_sc_hd__a32o_1 _4104_ (.A1(net272),
    .A2(_3424_),
    .A3(_3649_),
    .B1(_3670_),
    .B2(_3671_),
    .X(_3672_));
 sky130_fd_sc_hd__and3_1 _4105_ (.A(\mul_wb.lob_4.L[7] ),
    .B(_3383_),
    .C(_3399_),
    .X(_3673_));
 sky130_fd_sc_hd__a22o_1 _4106_ (.A1(\mul_wb.lob_4.L[4] ),
    .A2(net249),
    .B1(_3570_),
    .B2(\mul_wb.lob_4.L[5] ),
    .X(_3674_));
 sky130_fd_sc_hd__o21ai_1 _4107_ (.A1(_3673_),
    .A2(_3674_),
    .B1(_3424_),
    .Y(_3675_));
 sky130_fd_sc_hd__a32o_1 _4108_ (.A1(net268),
    .A2(_3412_),
    .A3(_3563_),
    .B1(_3565_),
    .B2(_3450_),
    .X(_3676_));
 sky130_fd_sc_hd__or4_1 _4109_ (.A(_3368_),
    .B(_3400_),
    .C(_3411_),
    .D(_3416_),
    .X(_3677_));
 sky130_fd_sc_hd__nand2_1 _4110_ (.A(\mul_wb.lob_4.L[8] ),
    .B(net246),
    .Y(_3678_));
 sky130_fd_sc_hd__or4_1 _4111_ (.A(_3369_),
    .B(net246),
    .C(_3405_),
    .D(_3409_),
    .X(_3679_));
 sky130_fd_sc_hd__a21o_1 _4112_ (.A1(_3678_),
    .A2(_3679_),
    .B1(_3445_),
    .X(_3680_));
 sky130_fd_sc_hd__or3_1 _4113_ (.A(_3370_),
    .B(_3456_),
    .C(_3576_),
    .X(_3681_));
 sky130_fd_sc_hd__a31o_1 _4114_ (.A1(_3677_),
    .A2(_3680_),
    .A3(_3681_),
    .B1(_3425_),
    .X(_3682_));
 sky130_fd_sc_hd__and4bb_4 _4115_ (.A_N(_3672_),
    .B_N(_3676_),
    .C(_3682_),
    .D(_3675_),
    .X(_3683_));
 sky130_fd_sc_hd__nor2_1 _4116_ (.A(net176),
    .B(net208),
    .Y(_3684_));
 sky130_fd_sc_hd__nand2_1 _4117_ (.A(_3666_),
    .B(_3684_),
    .Y(_3685_));
 sky130_fd_sc_hd__xnor2_2 _4118_ (.A(_3666_),
    .B(_3684_),
    .Y(_3686_));
 sky130_fd_sc_hd__or2_1 _4119_ (.A(_3614_),
    .B(net173),
    .X(_3687_));
 sky130_fd_sc_hd__and2_1 _4120_ (.A(net270),
    .B(_3526_),
    .X(_3688_));
 sky130_fd_sc_hd__a32o_1 _4121_ (.A1(net238),
    .A2(_3596_),
    .A3(_3688_),
    .B1(net243),
    .B2(\mul_wb.lob_4.L[6] ),
    .X(_3689_));
 sky130_fd_sc_hd__and4_1 _4122_ (.A(net273),
    .B(_3515_),
    .C(net239),
    .D(net238),
    .X(_3690_));
 sky130_fd_sc_hd__a221o_1 _4123_ (.A1(net275),
    .A2(_3626_),
    .B1(_3689_),
    .B2(_3542_),
    .C1(_3690_),
    .X(_3691_));
 sky130_fd_sc_hd__and2_1 _4124_ (.A(net274),
    .B(_3593_),
    .X(_3692_));
 sky130_fd_sc_hd__and3_1 _4125_ (.A(\mul_wb.lob_4.L[8] ),
    .B(_3488_),
    .C(net239),
    .X(_3693_));
 sky130_fd_sc_hd__a221o_1 _4126_ (.A1(net272),
    .A2(_3599_),
    .B1(_3600_),
    .B2(\mul_wb.lob_4.L[7] ),
    .C1(_3693_),
    .X(_3694_));
 sky130_fd_sc_hd__a22o_1 _4127_ (.A1(\mul_wb.lob_4.L[4] ),
    .A2(net245),
    .B1(_3589_),
    .B2(\mul_wb.lob_4.L[5] ),
    .X(_3695_));
 sky130_fd_sc_hd__a221o_1 _4128_ (.A1(\mul_wb.lob_4.L[9] ),
    .A2(_3592_),
    .B1(_3594_),
    .B2(_3531_),
    .C1(_3695_),
    .X(_3696_));
 sky130_fd_sc_hd__o41ai_4 _4129_ (.A1(_3691_),
    .A2(_3692_),
    .A3(_3694_),
    .A4(_3696_),
    .B1(_3521_),
    .Y(_3697_));
 sky130_fd_sc_hd__nor2_1 _4130_ (.A(net177),
    .B(net207),
    .Y(_3698_));
 sky130_fd_sc_hd__and2b_1 _4131_ (.A_N(_3687_),
    .B(_3698_),
    .X(_3699_));
 sky130_fd_sc_hd__xnor2_1 _4132_ (.A(_3687_),
    .B(_3698_),
    .Y(_3700_));
 sky130_fd_sc_hd__nand2_1 _4133_ (.A(_3659_),
    .B(_3700_),
    .Y(_3701_));
 sky130_fd_sc_hd__or2_1 _4134_ (.A(_3659_),
    .B(_3700_),
    .X(_3702_));
 sky130_fd_sc_hd__nand2_1 _4135_ (.A(_3701_),
    .B(_3702_),
    .Y(_3703_));
 sky130_fd_sc_hd__xor2_2 _4136_ (.A(_3686_),
    .B(_3703_),
    .X(_3704_));
 sky130_fd_sc_hd__nor2_1 _4137_ (.A(_3617_),
    .B(_3662_),
    .Y(_3705_));
 sky130_fd_sc_hd__xnor2_1 _4138_ (.A(_3704_),
    .B(_3705_),
    .Y(_3706_));
 sky130_fd_sc_hd__xnor2_1 _4139_ (.A(_3665_),
    .B(_3706_),
    .Y(\mul_wb.reg_p[3] ));
 sky130_fd_sc_hd__nor2_1 _4140_ (.A(net210),
    .B(net173),
    .Y(_3707_));
 sky130_fd_sc_hd__or4_1 _4141_ (.A(_3367_),
    .B(_3400_),
    .C(_3411_),
    .D(_3416_),
    .X(_3708_));
 sky130_fd_sc_hd__or3_1 _4142_ (.A(_3371_),
    .B(_3384_),
    .C(_3400_),
    .X(_3709_));
 sky130_fd_sc_hd__nand2_1 _4143_ (.A(\mul_wb.lob_4.L[9] ),
    .B(net246),
    .Y(_3710_));
 sky130_fd_sc_hd__or4_1 _4144_ (.A(_3368_),
    .B(net246),
    .C(_3405_),
    .D(_3409_),
    .X(_3711_));
 sky130_fd_sc_hd__a21o_1 _4145_ (.A1(_3710_),
    .A2(_3711_),
    .B1(_3445_),
    .X(_3712_));
 sky130_fd_sc_hd__nand2_1 _4146_ (.A(\mul_wb.lob_4.L[6] ),
    .B(_3570_),
    .Y(_3713_));
 sky130_fd_sc_hd__nand2_1 _4147_ (.A(\mul_wb.lob_4.L[5] ),
    .B(net249),
    .Y(_3714_));
 sky130_fd_sc_hd__or4_1 _4148_ (.A(_3366_),
    .B(_3418_),
    .C(_3445_),
    .D(_3447_),
    .X(_3715_));
 sky130_fd_sc_hd__or3_1 _4149_ (.A(_3369_),
    .B(_3456_),
    .C(_3576_),
    .X(_3716_));
 sky130_fd_sc_hd__a41o_1 _4150_ (.A1(_3708_),
    .A2(_3713_),
    .A3(_3714_),
    .A4(_3715_),
    .B1(_3431_),
    .X(_3717_));
 sky130_fd_sc_hd__a31o_1 _4151_ (.A1(_3709_),
    .A2(_3712_),
    .A3(_3716_),
    .B1(_3431_),
    .X(_3718_));
 sky130_fd_sc_hd__and2_1 _4152_ (.A(\mul_wb.lob_4.L[7] ),
    .B(net250),
    .X(_3719_));
 sky130_fd_sc_hd__a41o_1 _4153_ (.A1(net268),
    .A2(_3443_),
    .A3(_3446_),
    .A4(_3448_),
    .B1(_3719_),
    .X(_3720_));
 sky130_fd_sc_hd__a22oi_2 _4154_ (.A1(_3649_),
    .A2(_3669_),
    .B1(_3720_),
    .B2(_3573_),
    .Y(_3721_));
 sky130_fd_sc_hd__and3_4 _4155_ (.A(_3717_),
    .B(_3718_),
    .C(_3721_),
    .X(_3722_));
 sky130_fd_sc_hd__nor2_1 _4156_ (.A(net176),
    .B(net206),
    .Y(_3723_));
 sky130_fd_sc_hd__nand2_1 _4157_ (.A(_3707_),
    .B(_3723_),
    .Y(_3724_));
 sky130_fd_sc_hd__xnor2_1 _4158_ (.A(_3707_),
    .B(_3723_),
    .Y(_3725_));
 sky130_fd_sc_hd__and2_1 _4159_ (.A(net273),
    .B(_3593_),
    .X(_3726_));
 sky130_fd_sc_hd__and2_1 _4160_ (.A(\mul_wb.lob_4.L[10] ),
    .B(_3592_),
    .X(_3727_));
 sky130_fd_sc_hd__nor2_1 _4161_ (.A(_3370_),
    .B(_3489_),
    .Y(_3728_));
 sky130_fd_sc_hd__and2_1 _4162_ (.A(net274),
    .B(_3507_),
    .X(_3729_));
 sky130_fd_sc_hd__nand2_1 _4163_ (.A(net272),
    .B(_3515_),
    .Y(_3730_));
 sky130_fd_sc_hd__or3_1 _4164_ (.A(_3364_),
    .B(_3515_),
    .C(_3523_),
    .X(_3731_));
 sky130_fd_sc_hd__a21boi_1 _4165_ (.A1(_3730_),
    .A2(_3731_),
    .B1_N(_3529_),
    .Y(_3732_));
 sky130_fd_sc_hd__o21a_1 _4166_ (.A1(_3729_),
    .A2(_3732_),
    .B1(_3544_),
    .X(_3733_));
 sky130_fd_sc_hd__o21a_1 _4167_ (.A1(_3728_),
    .A2(_3733_),
    .B1(net239),
    .X(_3734_));
 sky130_fd_sc_hd__and3_1 _4168_ (.A(\mul_wb.lob_4.L[6] ),
    .B(net244),
    .C(_3495_),
    .X(_3735_));
 sky130_fd_sc_hd__a221o_1 _4169_ (.A1(\mul_wb.lob_4.L[5] ),
    .A2(net245),
    .B1(_3601_),
    .B2(\mul_wb.lob_4.L[7] ),
    .C1(_3735_),
    .X(_3736_));
 sky130_fd_sc_hd__a221o_1 _4170_ (.A1(net271),
    .A2(_3599_),
    .B1(_3600_),
    .B2(\mul_wb.lob_4.L[8] ),
    .C1(_3736_),
    .X(_3737_));
 sky130_fd_sc_hd__or4_4 _4171_ (.A(_3726_),
    .B(_3727_),
    .C(_3734_),
    .D(_3737_),
    .X(_3738_));
 sky130_fd_sc_hd__nand2_1 _4172_ (.A(_3526_),
    .B(_3738_),
    .Y(_3739_));
 sky130_fd_sc_hd__or3b_1 _4173_ (.A(net177),
    .B(_3527_),
    .C_N(_3738_),
    .X(_3740_));
 sky130_fd_sc_hd__a21oi_1 _4174_ (.A1(_3608_),
    .A2(_3613_),
    .B1(net208),
    .Y(_3741_));
 sky130_fd_sc_hd__a21oi_2 _4175_ (.A1(_3583_),
    .A2(_3586_),
    .B1(net207),
    .Y(_3742_));
 sky130_fd_sc_hd__nand2_1 _4176_ (.A(_3741_),
    .B(_3742_),
    .Y(_3743_));
 sky130_fd_sc_hd__xnor2_1 _4177_ (.A(_3741_),
    .B(_3742_),
    .Y(_3744_));
 sky130_fd_sc_hd__xnor2_1 _4178_ (.A(_3740_),
    .B(_3744_),
    .Y(_3745_));
 sky130_fd_sc_hd__nor2_1 _4179_ (.A(_3685_),
    .B(_3745_),
    .Y(_3746_));
 sky130_fd_sc_hd__xor2_1 _4180_ (.A(_3685_),
    .B(_3745_),
    .X(_3747_));
 sky130_fd_sc_hd__xnor2_1 _4181_ (.A(_3699_),
    .B(_3747_),
    .Y(_3748_));
 sky130_fd_sc_hd__nor2_1 _4182_ (.A(_3725_),
    .B(_3748_),
    .Y(_3749_));
 sky130_fd_sc_hd__xnor2_1 _4183_ (.A(_3725_),
    .B(_3748_),
    .Y(_3750_));
 sky130_fd_sc_hd__o21a_1 _4184_ (.A1(_3686_),
    .A2(_3703_),
    .B1(_3701_),
    .X(_3751_));
 sky130_fd_sc_hd__or2_1 _4185_ (.A(_3750_),
    .B(_3751_),
    .X(_3752_));
 sky130_fd_sc_hd__xor2_1 _4186_ (.A(_3750_),
    .B(_3751_),
    .X(_3753_));
 sky130_fd_sc_hd__nand3_1 _4187_ (.A(_3662_),
    .B(_3704_),
    .C(_3753_),
    .Y(_3754_));
 sky130_fd_sc_hd__a21o_1 _4188_ (.A1(_3662_),
    .A2(_3704_),
    .B1(_3753_),
    .X(_3755_));
 sky130_fd_sc_hd__and4_1 _4189_ (.A(_3617_),
    .B(_3661_),
    .C(_3704_),
    .D(_3753_),
    .X(_3756_));
 sky130_fd_sc_hd__inv_2 _4190_ (.A(_3756_),
    .Y(_3757_));
 sky130_fd_sc_hd__a32o_1 _4191_ (.A1(_3617_),
    .A2(_3661_),
    .A3(_3704_),
    .B1(_3754_),
    .B2(_3755_),
    .X(_3758_));
 sky130_fd_sc_hd__nand2_1 _4192_ (.A(_3757_),
    .B(_3758_),
    .Y(_3759_));
 sky130_fd_sc_hd__nor2_1 _4193_ (.A(_3664_),
    .B(_3706_),
    .Y(_3760_));
 sky130_fd_sc_hd__nor2_1 _4194_ (.A(_3620_),
    .B(_3760_),
    .Y(_3761_));
 sky130_fd_sc_hd__xnor2_1 _4195_ (.A(_3759_),
    .B(_3761_),
    .Y(\mul_wb.reg_p[4] ));
 sky130_fd_sc_hd__and2_1 _4196_ (.A(_3759_),
    .B(_3760_),
    .X(_3762_));
 sky130_fd_sc_hd__nor2_1 _4197_ (.A(_3620_),
    .B(_3762_),
    .Y(_3763_));
 sky130_fd_sc_hd__and4_1 _4198_ (.A(net273),
    .B(_3407_),
    .C(_3408_),
    .D(net241),
    .X(_3764_));
 sky130_fd_sc_hd__a221o_1 _4199_ (.A1(net270),
    .A2(_3565_),
    .B1(_3577_),
    .B2(net274),
    .C1(_3764_),
    .X(_3765_));
 sky130_fd_sc_hd__and2_1 _4200_ (.A(net272),
    .B(_3578_),
    .X(_3766_));
 sky130_fd_sc_hd__and4_1 _4201_ (.A(net268),
    .B(_3399_),
    .C(_3410_),
    .D(_3419_),
    .X(_3767_));
 sky130_fd_sc_hd__and3_1 _4202_ (.A(\mul_wb.lob_4.L[9] ),
    .B(_3383_),
    .C(_3399_),
    .X(_3768_));
 sky130_fd_sc_hd__and3_1 _4203_ (.A(net275),
    .B(net246),
    .C(net241),
    .X(_3769_));
 sky130_fd_sc_hd__and3_1 _4204_ (.A(\mul_wb.lob_4.L[7] ),
    .B(_3388_),
    .C(_3396_),
    .X(_3770_));
 sky130_fd_sc_hd__a221o_1 _4205_ (.A1(\mul_wb.lob_4.L[6] ),
    .A2(net248),
    .B1(_3568_),
    .B2(\mul_wb.lob_4.L[8] ),
    .C1(_3770_),
    .X(_3771_));
 sky130_fd_sc_hd__or4_1 _4206_ (.A(_3767_),
    .B(_3768_),
    .C(_3769_),
    .D(_3771_),
    .X(_3772_));
 sky130_fd_sc_hd__o31ai_2 _4207_ (.A1(_3765_),
    .A2(_3766_),
    .A3(_3772_),
    .B1(_3429_),
    .Y(_3773_));
 sky130_fd_sc_hd__nor2_1 _4208_ (.A(net175),
    .B(net204),
    .Y(_3774_));
 sky130_fd_sc_hd__or2_1 _4209_ (.A(net210),
    .B(net208),
    .X(_3775_));
 sky130_fd_sc_hd__a32o_1 _4210_ (.A1(net275),
    .A2(_3488_),
    .A3(_3502_),
    .B1(net243),
    .B2(\mul_wb.lob_4.L[8] ),
    .X(_3776_));
 sky130_fd_sc_hd__a22o_1 _4211_ (.A1(\mul_wb.lob_4.L[6] ),
    .A2(net245),
    .B1(_3589_),
    .B2(\mul_wb.lob_4.L[7] ),
    .X(_3777_));
 sky130_fd_sc_hd__a221o_1 _4212_ (.A1(\mul_wb.lob_4.L[9] ),
    .A2(_3600_),
    .B1(_3776_),
    .B2(_3542_),
    .C1(_3777_),
    .X(_3778_));
 sky130_fd_sc_hd__a22o_1 _4213_ (.A1(net270),
    .A2(_3590_),
    .B1(_3626_),
    .B2(net273),
    .X(_3779_));
 sky130_fd_sc_hd__nor3_1 _4214_ (.A(_3364_),
    .B(_3511_),
    .C(_3515_),
    .Y(_3780_));
 sky130_fd_sc_hd__a21o_1 _4215_ (.A1(net272),
    .A2(_3511_),
    .B1(_3780_),
    .X(_3781_));
 sky130_fd_sc_hd__a32o_1 _4216_ (.A1(_3508_),
    .A2(_3514_),
    .A3(_3781_),
    .B1(_3592_),
    .B2(net274),
    .X(_3782_));
 sky130_fd_sc_hd__o31ai_4 _4217_ (.A1(_3778_),
    .A2(_3779_),
    .A3(_3782_),
    .B1(_3523_),
    .Y(_3783_));
 sky130_fd_sc_hd__o21ai_1 _4218_ (.A1(net177),
    .A2(net202),
    .B1(_3775_),
    .Y(_3784_));
 sky130_fd_sc_hd__or3_1 _4219_ (.A(net177),
    .B(_3775_),
    .C(net202),
    .X(_3785_));
 sky130_fd_sc_hd__and2_1 _4220_ (.A(_3784_),
    .B(_3785_),
    .X(_3786_));
 sky130_fd_sc_hd__xnor2_1 _4221_ (.A(_3774_),
    .B(_3786_),
    .Y(_3787_));
 sky130_fd_sc_hd__o21ai_1 _4222_ (.A1(_3740_),
    .A2(_3744_),
    .B1(_3743_),
    .Y(_3788_));
 sky130_fd_sc_hd__or3b_1 _4223_ (.A(_3527_),
    .B(net174),
    .C_N(_3738_),
    .X(_3789_));
 sky130_fd_sc_hd__a21o_1 _4224_ (.A1(_3648_),
    .A2(_3656_),
    .B1(net207),
    .X(_3790_));
 sky130_fd_sc_hd__a21oi_1 _4225_ (.A1(_3608_),
    .A2(_3613_),
    .B1(net206),
    .Y(_0241_));
 sky130_fd_sc_hd__xnor2_1 _4226_ (.A(_3790_),
    .B(_0241_),
    .Y(_0242_));
 sky130_fd_sc_hd__nand2b_1 _4227_ (.A_N(_3789_),
    .B(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hd__xnor2_1 _4228_ (.A(_3789_),
    .B(_0242_),
    .Y(_0244_));
 sky130_fd_sc_hd__and3_1 _4229_ (.A(_3707_),
    .B(_3723_),
    .C(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__xnor2_1 _4230_ (.A(_3724_),
    .B(_0244_),
    .Y(_0246_));
 sky130_fd_sc_hd__and2_1 _4231_ (.A(_3788_),
    .B(_0246_),
    .X(_0247_));
 sky130_fd_sc_hd__xor2_1 _4232_ (.A(_3788_),
    .B(_0246_),
    .X(_0248_));
 sky130_fd_sc_hd__nand2b_1 _4233_ (.A_N(_3787_),
    .B(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__xnor2_1 _4234_ (.A(_3787_),
    .B(_0248_),
    .Y(_0250_));
 sky130_fd_sc_hd__and2_1 _4235_ (.A(_3749_),
    .B(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__or2_1 _4236_ (.A(_3749_),
    .B(_0250_),
    .X(_0252_));
 sky130_fd_sc_hd__xor2_1 _4237_ (.A(_3749_),
    .B(_0250_),
    .X(_0253_));
 sky130_fd_sc_hd__a21o_1 _4238_ (.A1(_3699_),
    .A2(_3747_),
    .B1(_3746_),
    .X(_0254_));
 sky130_fd_sc_hd__xnor2_2 _4239_ (.A(_0253_),
    .B(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__and3_1 _4240_ (.A(_3752_),
    .B(_3754_),
    .C(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__nor2_1 _4241_ (.A(_3754_),
    .B(_0255_),
    .Y(_0257_));
 sky130_fd_sc_hd__or2_1 _4242_ (.A(_3754_),
    .B(_0255_),
    .X(_0258_));
 sky130_fd_sc_hd__nor2_1 _4243_ (.A(_3752_),
    .B(_0255_),
    .Y(_0259_));
 sky130_fd_sc_hd__or2_1 _4244_ (.A(_0256_),
    .B(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__or2_1 _4245_ (.A(_0257_),
    .B(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__or2_1 _4246_ (.A(_3757_),
    .B(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__xnor2_1 _4247_ (.A(_3757_),
    .B(_0261_),
    .Y(_0263_));
 sky130_fd_sc_hd__xnor2_1 _4248_ (.A(_3763_),
    .B(_0263_),
    .Y(\mul_wb.reg_p[5] ));
 sky130_fd_sc_hd__a32o_1 _4249_ (.A1(net269),
    .A2(_3543_),
    .A3(net238),
    .B1(\mul_wb.lob_4.L[7] ),
    .B2(net245),
    .X(_0264_));
 sky130_fd_sc_hd__a221o_1 _4250_ (.A1(\mul_wb.lob_4.L[12] ),
    .A2(_3592_),
    .B1(_3626_),
    .B2(net272),
    .C1(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__and2_1 _4251_ (.A(net270),
    .B(_3593_),
    .X(_0266_));
 sky130_fd_sc_hd__or4_1 _4252_ (.A(_3368_),
    .B(_3487_),
    .C(_3489_),
    .D(net243),
    .X(_0267_));
 sky130_fd_sc_hd__nand2_1 _4253_ (.A(\mul_wb.lob_4.L[9] ),
    .B(_3493_),
    .Y(_0268_));
 sky130_fd_sc_hd__a21oi_1 _4254_ (.A1(_0267_),
    .A2(_0268_),
    .B1(_3495_),
    .Y(_0269_));
 sky130_fd_sc_hd__a22o_1 _4255_ (.A1(\mul_wb.lob_4.L[8] ),
    .A2(_3495_),
    .B1(_3632_),
    .B2(\mul_wb.lob_4.L[10] ),
    .X(_0270_));
 sky130_fd_sc_hd__o21a_1 _4256_ (.A1(_0269_),
    .A2(_0270_),
    .B1(net244),
    .X(_0271_));
 sky130_fd_sc_hd__o31ai_2 _4257_ (.A1(_0265_),
    .A2(_0266_),
    .A3(_0271_),
    .B1(_3515_),
    .Y(_0272_));
 sky130_fd_sc_hd__nor2_1 _4258_ (.A(net177),
    .B(net200),
    .Y(_0273_));
 sky130_fd_sc_hd__o21a_1 _4259_ (.A1(_0245_),
    .A2(_0247_),
    .B1(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__nor3_1 _4260_ (.A(_0245_),
    .B(_0247_),
    .C(_0273_),
    .Y(_0275_));
 sky130_fd_sc_hd__nor2_1 _4261_ (.A(_0274_),
    .B(_0275_),
    .Y(_0276_));
 sky130_fd_sc_hd__nand2_1 _4262_ (.A(\mul_wb.lob_4.L[9] ),
    .B(net250),
    .Y(_0277_));
 sky130_fd_sc_hd__a2111o_1 _4263_ (.A1(_3381_),
    .A2(_3382_),
    .B1(net250),
    .C1(_3402_),
    .D1(_3368_),
    .X(_0278_));
 sky130_fd_sc_hd__a21oi_1 _4264_ (.A1(_0277_),
    .A2(_0278_),
    .B1(_3388_),
    .Y(_0279_));
 sky130_fd_sc_hd__a32o_1 _4265_ (.A1(net275),
    .A2(_3383_),
    .A3(_3391_),
    .B1(_3388_),
    .B2(\mul_wb.lob_4.L[8] ),
    .X(_0280_));
 sky130_fd_sc_hd__o21a_1 _4266_ (.A1(_0279_),
    .A2(_0280_),
    .B1(_3396_),
    .X(_0281_));
 sky130_fd_sc_hd__and4_1 _4267_ (.A(net270),
    .B(_3399_),
    .C(_3410_),
    .D(_3415_),
    .X(_0282_));
 sky130_fd_sc_hd__and4_1 _4268_ (.A(net272),
    .B(_3407_),
    .C(_3408_),
    .D(net241),
    .X(_0283_));
 sky130_fd_sc_hd__a32o_1 _4269_ (.A1(net268),
    .A2(net241),
    .A3(_3446_),
    .B1(\mul_wb.lob_4.L[7] ),
    .B2(net248),
    .X(_0284_));
 sky130_fd_sc_hd__a2111o_1 _4270_ (.A1(net273),
    .A2(_3577_),
    .B1(_0282_),
    .C1(_0283_),
    .D1(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__o21ai_1 _4271_ (.A1(_0281_),
    .A2(_0285_),
    .B1(_3417_),
    .Y(_0286_));
 sky130_fd_sc_hd__nor2_2 _4272_ (.A(net175),
    .B(net198),
    .Y(_0287_));
 sky130_fd_sc_hd__nor2_1 _4273_ (.A(net209),
    .B(net206),
    .Y(_0288_));
 sky130_fd_sc_hd__o21bai_2 _4274_ (.A1(net174),
    .A2(net202),
    .B1_N(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__or3b_1 _4275_ (.A(net174),
    .B(net202),
    .C_N(_0288_),
    .X(_0290_));
 sky130_fd_sc_hd__nand2_1 _4276_ (.A(_0289_),
    .B(_0290_),
    .Y(_0291_));
 sky130_fd_sc_hd__xnor2_2 _4277_ (.A(_0287_),
    .B(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__o31ai_4 _4278_ (.A1(_3614_),
    .A2(net206),
    .A3(_3790_),
    .B1(_0243_),
    .Y(_0293_));
 sky130_fd_sc_hd__a21bo_1 _4279_ (.A1(_3774_),
    .A2(_3784_),
    .B1_N(_3785_),
    .X(_0294_));
 sky130_fd_sc_hd__or3b_2 _4280_ (.A(_3527_),
    .B(net173),
    .C_N(_3738_),
    .X(_0295_));
 sky130_fd_sc_hd__or2_2 _4281_ (.A(net208),
    .B(net207),
    .X(_0296_));
 sky130_fd_sc_hd__a21oi_1 _4282_ (.A1(_3608_),
    .A2(_3613_),
    .B1(net204),
    .Y(_0297_));
 sky130_fd_sc_hd__xnor2_2 _4283_ (.A(_0296_),
    .B(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__nand2b_1 _4284_ (.A_N(_0295_),
    .B(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__xor2_2 _4285_ (.A(_0295_),
    .B(_0298_),
    .X(_0300_));
 sky130_fd_sc_hd__and2b_1 _4286_ (.A_N(_0300_),
    .B(_0294_),
    .X(_0301_));
 sky130_fd_sc_hd__xnor2_2 _4287_ (.A(_0294_),
    .B(_0300_),
    .Y(_0302_));
 sky130_fd_sc_hd__and2_1 _4288_ (.A(_0293_),
    .B(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__xor2_2 _4289_ (.A(_0293_),
    .B(_0302_),
    .X(_0304_));
 sky130_fd_sc_hd__nand2_1 _4290_ (.A(_0292_),
    .B(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__xor2_2 _4291_ (.A(_0292_),
    .B(_0304_),
    .X(_0306_));
 sky130_fd_sc_hd__and2b_1 _4292_ (.A_N(_0249_),
    .B(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__xnor2_2 _4293_ (.A(_0249_),
    .B(_0306_),
    .Y(_0308_));
 sky130_fd_sc_hd__xor2_2 _4294_ (.A(_0276_),
    .B(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__a21oi_2 _4295_ (.A1(_0252_),
    .A2(_0254_),
    .B1(_0251_),
    .Y(_0310_));
 sky130_fd_sc_hd__and2b_1 _4296_ (.A_N(_0310_),
    .B(_0309_),
    .X(_0311_));
 sky130_fd_sc_hd__xnor2_2 _4297_ (.A(_0309_),
    .B(_0310_),
    .Y(_0312_));
 sky130_fd_sc_hd__nand2_1 _4298_ (.A(_0259_),
    .B(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__xnor2_1 _4299_ (.A(_0259_),
    .B(_0312_),
    .Y(_0314_));
 sky130_fd_sc_hd__or2_1 _4300_ (.A(_0258_),
    .B(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__nand2_1 _4301_ (.A(_0258_),
    .B(_0314_),
    .Y(_0316_));
 sky130_fd_sc_hd__nand2_1 _4302_ (.A(_0315_),
    .B(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__or4_1 _4303_ (.A(_3757_),
    .B(_0257_),
    .C(_0260_),
    .D(_0314_),
    .X(_0318_));
 sky130_fd_sc_hd__xnor2_1 _4304_ (.A(_0262_),
    .B(_0317_),
    .Y(_0319_));
 sky130_fd_sc_hd__and2_1 _4305_ (.A(_3762_),
    .B(_0263_),
    .X(_0320_));
 sky130_fd_sc_hd__nor2_1 _4306_ (.A(_3620_),
    .B(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__xnor2_1 _4307_ (.A(_0319_),
    .B(_0321_),
    .Y(\mul_wb.reg_p[6] ));
 sky130_fd_sc_hd__nand2_1 _4308_ (.A(_0319_),
    .B(_0320_),
    .Y(_0322_));
 sky130_fd_sc_hd__nand2_1 _4309_ (.A(net252),
    .B(_0322_),
    .Y(_0323_));
 sky130_fd_sc_hd__or2_1 _4310_ (.A(net174),
    .B(net200),
    .X(_0324_));
 sky130_fd_sc_hd__a32o_1 _4311_ (.A1(net271),
    .A2(_3507_),
    .A3(_3544_),
    .B1(\mul_wb.lob_4.L[12] ),
    .B2(_3488_),
    .X(_0325_));
 sky130_fd_sc_hd__nor2_1 _4312_ (.A(_3371_),
    .B(net244),
    .Y(_0326_));
 sky130_fd_sc_hd__a221o_1 _4313_ (.A1(\mul_wb.lob_4.L[7] ),
    .A2(_3498_),
    .B1(_3601_),
    .B2(\mul_wb.lob_4.L[10] ),
    .C1(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__a21o_1 _4314_ (.A1(net239),
    .A2(_0325_),
    .B1(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__and4_1 _4315_ (.A(net268),
    .B(_3503_),
    .C(_3508_),
    .D(_3513_),
    .X(_0329_));
 sky130_fd_sc_hd__a22o_1 _4316_ (.A1(\mul_wb.lob_4.L[9] ),
    .A2(_3495_),
    .B1(_3632_),
    .B2(net274),
    .X(_0330_));
 sky130_fd_sc_hd__a221o_1 _4317_ (.A1(net272),
    .A2(_3592_),
    .B1(_0330_),
    .B2(_3513_),
    .C1(_0329_),
    .X(_0331_));
 sky130_fd_sc_hd__o21ai_2 _4318_ (.A1(_0328_),
    .A2(_0331_),
    .B1(_3511_),
    .Y(_0332_));
 sky130_fd_sc_hd__or3_1 _4319_ (.A(net177),
    .B(_0324_),
    .C(net196),
    .X(_0333_));
 sky130_fd_sc_hd__o21ai_1 _4320_ (.A1(net177),
    .A2(net196),
    .B1(_0324_),
    .Y(_0334_));
 sky130_fd_sc_hd__and2_1 _4321_ (.A(_0333_),
    .B(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__o21a_2 _4322_ (.A1(_0301_),
    .A2(_0303_),
    .B1(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__nor3_1 _4323_ (.A(_0301_),
    .B(_0303_),
    .C(_0335_),
    .Y(_0337_));
 sky130_fd_sc_hd__nor2_1 _4324_ (.A(_0336_),
    .B(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__a32o_1 _4325_ (.A1(net274),
    .A2(_3383_),
    .A3(_3391_),
    .B1(_3388_),
    .B2(\mul_wb.lob_4.L[9] ),
    .X(_0339_));
 sky130_fd_sc_hd__and4_1 _4326_ (.A(net270),
    .B(_3407_),
    .C(_3408_),
    .D(_3444_),
    .X(_0340_));
 sky130_fd_sc_hd__a221o_2 _4327_ (.A1(\mul_wb.lob_4.L[13] ),
    .A2(_3577_),
    .B1(_0339_),
    .B2(_3398_),
    .C1(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__and2_1 _4328_ (.A(net275),
    .B(_3568_),
    .X(_0342_));
 sky130_fd_sc_hd__a22o_1 _4329_ (.A1(\mul_wb.lob_4.L[8] ),
    .A2(net248),
    .B1(net247),
    .B2(\mul_wb.lob_4.L[7] ),
    .X(_0343_));
 sky130_fd_sc_hd__a31o_1 _4330_ (.A1(\mul_wb.lob_4.L[12] ),
    .A2(_3401_),
    .A3(_3444_),
    .B1(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__a211o_2 _4331_ (.A1(net268),
    .A2(_3412_),
    .B1(_0342_),
    .C1(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__o21ai_4 _4332_ (.A1(_0341_),
    .A2(_0345_),
    .B1(_3415_),
    .Y(_0346_));
 sky130_fd_sc_hd__nor2_2 _4333_ (.A(net175),
    .B(net195),
    .Y(_0347_));
 sky130_fd_sc_hd__or2_1 _4334_ (.A(net209),
    .B(net204),
    .X(_0348_));
 sky130_fd_sc_hd__o21ai_2 _4335_ (.A1(net173),
    .A2(net202),
    .B1(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__or3_1 _4336_ (.A(net173),
    .B(net202),
    .C(_0348_),
    .X(_0350_));
 sky130_fd_sc_hd__nand2_2 _4337_ (.A(_0349_),
    .B(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__xnor2_4 _4338_ (.A(_0347_),
    .B(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__o31ai_4 _4339_ (.A1(_3614_),
    .A2(net204),
    .A3(_0296_),
    .B1(_0299_),
    .Y(_0353_));
 sky130_fd_sc_hd__a21boi_4 _4340_ (.A1(_0287_),
    .A2(_0289_),
    .B1_N(_0290_),
    .Y(_0354_));
 sky130_fd_sc_hd__and3b_2 _4341_ (.A_N(net208),
    .B(_3738_),
    .C(_3526_),
    .X(_0355_));
 sky130_fd_sc_hd__nor2_2 _4342_ (.A(net207),
    .B(net206),
    .Y(_0356_));
 sky130_fd_sc_hd__a21oi_2 _4343_ (.A1(_3608_),
    .A2(_3613_),
    .B1(net198),
    .Y(_0357_));
 sky130_fd_sc_hd__xor2_4 _4344_ (.A(_0356_),
    .B(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__xnor2_4 _4345_ (.A(_0355_),
    .B(_0358_),
    .Y(_0359_));
 sky130_fd_sc_hd__nor2_1 _4346_ (.A(_0354_),
    .B(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hd__xor2_4 _4347_ (.A(_0354_),
    .B(_0359_),
    .X(_0361_));
 sky130_fd_sc_hd__xor2_4 _4348_ (.A(_0353_),
    .B(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__nand2_1 _4349_ (.A(_0352_),
    .B(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__xor2_2 _4350_ (.A(_0352_),
    .B(_0362_),
    .X(_0364_));
 sky130_fd_sc_hd__xnor2_2 _4351_ (.A(_0305_),
    .B(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__xnor2_2 _4352_ (.A(_0338_),
    .B(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__a21oi_2 _4353_ (.A1(_0276_),
    .A2(_0308_),
    .B1(_0307_),
    .Y(_0367_));
 sky130_fd_sc_hd__nor2_1 _4354_ (.A(_0366_),
    .B(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__xor2_2 _4355_ (.A(_0366_),
    .B(_0367_),
    .X(_0369_));
 sky130_fd_sc_hd__xnor2_2 _4356_ (.A(_0274_),
    .B(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__a21oi_1 _4357_ (.A1(_0259_),
    .A2(_0312_),
    .B1(_0311_),
    .Y(_0371_));
 sky130_fd_sc_hd__xnor2_1 _4358_ (.A(_0370_),
    .B(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__a21o_1 _4359_ (.A1(_0315_),
    .A2(_0318_),
    .B1(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__nand3_1 _4360_ (.A(_0315_),
    .B(_0318_),
    .C(_0372_),
    .Y(_0374_));
 sky130_fd_sc_hd__and2_1 _4361_ (.A(_0373_),
    .B(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__xnor2_1 _4362_ (.A(_0323_),
    .B(_0375_),
    .Y(\mul_wb.reg_p[7] ));
 sky130_fd_sc_hd__nor3b_2 _4363_ (.A(_0310_),
    .B(_0370_),
    .C_N(_0309_),
    .Y(_0376_));
 sky130_fd_sc_hd__a21oi_2 _4364_ (.A1(_0274_),
    .A2(_0369_),
    .B1(_0368_),
    .Y(_0377_));
 sky130_fd_sc_hd__a21o_1 _4365_ (.A1(_0353_),
    .A2(_0361_),
    .B1(_0360_),
    .X(_0378_));
 sky130_fd_sc_hd__or4_4 _4366_ (.A(net174),
    .B(net173),
    .C(net200),
    .D(net196),
    .X(_0379_));
 sky130_fd_sc_hd__and2b_1 _4367_ (.A_N(_0379_),
    .B(_0333_),
    .X(_0380_));
 sky130_fd_sc_hd__and2b_2 _4368_ (.A_N(_0333_),
    .B(_0379_),
    .X(_0381_));
 sky130_fd_sc_hd__o22a_1 _4369_ (.A1(net173),
    .A2(net200),
    .B1(net196),
    .B2(net174),
    .X(_0382_));
 sky130_fd_sc_hd__or3_1 _4370_ (.A(_0380_),
    .B(_0381_),
    .C(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__and2b_1 _4371_ (.A_N(_0383_),
    .B(_0378_),
    .X(_0384_));
 sky130_fd_sc_hd__xnor2_2 _4372_ (.A(_0378_),
    .B(_0383_),
    .Y(_0385_));
 sky130_fd_sc_hd__a21o_1 _4373_ (.A1(net272),
    .A2(_3488_),
    .B1(_3636_),
    .X(_0386_));
 sky130_fd_sc_hd__nor2_1 _4374_ (.A(_3370_),
    .B(net244),
    .Y(_0387_));
 sky130_fd_sc_hd__a221o_1 _4375_ (.A1(net273),
    .A2(_3600_),
    .B1(_0386_),
    .B2(net239),
    .C1(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__a22o_1 _4376_ (.A1(net275),
    .A2(_3495_),
    .B1(_3499_),
    .B2(\mul_wb.lob_4.L[11] ),
    .X(_0389_));
 sky130_fd_sc_hd__a22o_1 _4377_ (.A1(net270),
    .A2(_3592_),
    .B1(_0389_),
    .B2(net244),
    .X(_0390_));
 sky130_fd_sc_hd__o21ai_2 _4378_ (.A1(_0388_),
    .A2(_0390_),
    .B1(_3507_),
    .Y(_0391_));
 sky130_fd_sc_hd__nor2_1 _4379_ (.A(_3475_),
    .B(net194),
    .Y(_0392_));
 sky130_fd_sc_hd__nand2_1 _4380_ (.A(net273),
    .B(_3567_),
    .Y(_0393_));
 sky130_fd_sc_hd__a22o_1 _4381_ (.A1(\mul_wb.lob_4.L[13] ),
    .A2(net246),
    .B1(_3407_),
    .B2(net268),
    .X(_0394_));
 sky130_fd_sc_hd__o2bb2a_1 _4382_ (.A1_N(_3444_),
    .A2_N(_0394_),
    .B1(_3370_),
    .B2(_3396_),
    .X(_0395_));
 sky130_fd_sc_hd__and3_1 _4383_ (.A(\mul_wb.lob_4.L[11] ),
    .B(_3389_),
    .C(_3390_),
    .X(_0396_));
 sky130_fd_sc_hd__a21oi_1 _4384_ (.A1(net275),
    .A2(_3388_),
    .B1(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__o2bb2a_1 _4385_ (.A1_N(net271),
    .A2_N(_3577_),
    .B1(_0397_),
    .B2(net249),
    .X(_0398_));
 sky130_fd_sc_hd__a31o_1 _4386_ (.A1(_0393_),
    .A2(_0395_),
    .A3(_0398_),
    .B1(_3409_),
    .X(_0399_));
 sky130_fd_sc_hd__nor2_1 _4387_ (.A(net175),
    .B(net192),
    .Y(_0400_));
 sky130_fd_sc_hd__o22a_1 _4388_ (.A1(net208),
    .A2(net202),
    .B1(net198),
    .B2(net209),
    .X(_0401_));
 sky130_fd_sc_hd__or4_1 _4389_ (.A(net209),
    .B(net208),
    .C(net202),
    .D(net198),
    .X(_0402_));
 sky130_fd_sc_hd__nand2b_1 _4390_ (.A_N(_0401_),
    .B(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__xnor2_1 _4391_ (.A(_0400_),
    .B(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__nand2_1 _4392_ (.A(_0392_),
    .B(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__or2_1 _4393_ (.A(_0392_),
    .B(_0404_),
    .X(_0406_));
 sky130_fd_sc_hd__and2_2 _4394_ (.A(_0405_),
    .B(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__a22o_2 _4395_ (.A1(_0356_),
    .A2(_0357_),
    .B1(_0358_),
    .B2(_0355_),
    .X(_0408_));
 sky130_fd_sc_hd__a21boi_4 _4396_ (.A1(_0347_),
    .A2(_0349_),
    .B1_N(_0350_),
    .Y(_0409_));
 sky130_fd_sc_hd__and3b_2 _4397_ (.A_N(net206),
    .B(_3738_),
    .C(_3526_),
    .X(_0410_));
 sky130_fd_sc_hd__or2_2 _4398_ (.A(net207),
    .B(net204),
    .X(_0411_));
 sky130_fd_sc_hd__a21oi_2 _4399_ (.A1(net212),
    .A2(net211),
    .B1(net195),
    .Y(_0412_));
 sky130_fd_sc_hd__or3_1 _4400_ (.A(_3614_),
    .B(net195),
    .C(_0411_),
    .X(_0413_));
 sky130_fd_sc_hd__xnor2_4 _4401_ (.A(_0411_),
    .B(_0412_),
    .Y(_0414_));
 sky130_fd_sc_hd__xnor2_4 _4402_ (.A(_0410_),
    .B(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__nor2_1 _4403_ (.A(_0409_),
    .B(_0415_),
    .Y(_0416_));
 sky130_fd_sc_hd__xor2_4 _4404_ (.A(_0409_),
    .B(_0415_),
    .X(_0417_));
 sky130_fd_sc_hd__xor2_4 _4405_ (.A(_0408_),
    .B(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__nand2_2 _4406_ (.A(_0407_),
    .B(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__xor2_4 _4407_ (.A(_0407_),
    .B(_0418_),
    .X(_0420_));
 sky130_fd_sc_hd__xnor2_2 _4408_ (.A(_0363_),
    .B(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__xnor2_2 _4409_ (.A(_0385_),
    .B(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__a32o_1 _4410_ (.A1(_0292_),
    .A2(_0304_),
    .A3(_0364_),
    .B1(_0365_),
    .B2(_0338_),
    .X(_0423_));
 sky130_fd_sc_hd__nand2b_1 _4411_ (.A_N(_0422_),
    .B(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__xnor2_2 _4412_ (.A(_0422_),
    .B(_0423_),
    .Y(_0425_));
 sky130_fd_sc_hd__xnor2_2 _4413_ (.A(_0336_),
    .B(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__or2_1 _4414_ (.A(_0377_),
    .B(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__xor2_2 _4415_ (.A(_0377_),
    .B(_0426_),
    .X(_0428_));
 sky130_fd_sc_hd__nand2_1 _4416_ (.A(_0376_),
    .B(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__xnor2_2 _4417_ (.A(_0376_),
    .B(_0428_),
    .Y(_0430_));
 sky130_fd_sc_hd__nor2_1 _4418_ (.A(_0313_),
    .B(_0370_),
    .Y(_0431_));
 sky130_fd_sc_hd__inv_2 _4419_ (.A(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__nand2_1 _4420_ (.A(_0373_),
    .B(_0432_),
    .Y(_0433_));
 sky130_fd_sc_hd__a21o_1 _4421_ (.A1(_0373_),
    .A2(_0432_),
    .B1(_0430_),
    .X(_0434_));
 sky130_fd_sc_hd__xnor2_2 _4422_ (.A(_0430_),
    .B(_0433_),
    .Y(_0435_));
 sky130_fd_sc_hd__o21a_1 _4423_ (.A1(_0322_),
    .A2(_0375_),
    .B1(net252),
    .X(_0436_));
 sky130_fd_sc_hd__xor2_1 _4424_ (.A(_0435_),
    .B(_0436_),
    .X(\mul_wb.reg_p[8] ));
 sky130_fd_sc_hd__a21oi_4 _4425_ (.A1(_0408_),
    .A2(_0417_),
    .B1(_0416_),
    .Y(_0437_));
 sky130_fd_sc_hd__a22o_1 _4426_ (.A1(net274),
    .A2(_3495_),
    .B1(_3632_),
    .B2(\mul_wb.lob_4.L[13] ),
    .X(_0438_));
 sky130_fd_sc_hd__and2_1 _4427_ (.A(_3513_),
    .B(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__a32o_1 _4428_ (.A1(net271),
    .A2(_3488_),
    .A3(_3502_),
    .B1(_3493_),
    .B2(net273),
    .X(_0440_));
 sky130_fd_sc_hd__a221o_1 _4429_ (.A1(net275),
    .A2(net245),
    .B1(_3542_),
    .B2(_0440_),
    .C1(_3594_),
    .X(_0441_));
 sky130_fd_sc_hd__o21ai_4 _4430_ (.A1(_0439_),
    .A2(_0441_),
    .B1(_3506_),
    .Y(_0442_));
 sky130_fd_sc_hd__nor2_2 _4431_ (.A(net177),
    .B(net191),
    .Y(_0443_));
 sky130_fd_sc_hd__o22a_1 _4432_ (.A1(net208),
    .A2(net200),
    .B1(net196),
    .B2(net173),
    .X(_0444_));
 sky130_fd_sc_hd__o22ai_1 _4433_ (.A1(net208),
    .A2(net200),
    .B1(net196),
    .B2(net173),
    .Y(_0445_));
 sky130_fd_sc_hd__nor4_1 _4434_ (.A(net173),
    .B(_3683_),
    .C(net200),
    .D(net196),
    .Y(_0446_));
 sky130_fd_sc_hd__nor2_2 _4435_ (.A(_0444_),
    .B(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__xor2_4 _4436_ (.A(_0443_),
    .B(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__nand2b_1 _4437_ (.A_N(_0379_),
    .B(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__xnor2_4 _4438_ (.A(_0379_),
    .B(_0448_),
    .Y(_0450_));
 sky130_fd_sc_hd__and2b_1 _4439_ (.A_N(_0437_),
    .B(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__xnor2_4 _4440_ (.A(_0437_),
    .B(_0450_),
    .Y(_0452_));
 sky130_fd_sc_hd__xor2_4 _4441_ (.A(_0381_),
    .B(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__a21bo_2 _4442_ (.A1(_0410_),
    .A2(_0414_),
    .B1_N(_0413_),
    .X(_0454_));
 sky130_fd_sc_hd__o31a_2 _4443_ (.A1(net175),
    .A2(net192),
    .A3(_0401_),
    .B1(_0402_),
    .X(_0455_));
 sky130_fd_sc_hd__or3b_4 _4444_ (.A(_3527_),
    .B(net204),
    .C_N(_3738_),
    .X(_0456_));
 sky130_fd_sc_hd__nor2_2 _4445_ (.A(net207),
    .B(net198),
    .Y(_0457_));
 sky130_fd_sc_hd__a21oi_2 _4446_ (.A1(net212),
    .A2(net211),
    .B1(net192),
    .Y(_0458_));
 sky130_fd_sc_hd__nand2_1 _4447_ (.A(_0457_),
    .B(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__xnor2_4 _4448_ (.A(_0457_),
    .B(_0458_),
    .Y(_0460_));
 sky130_fd_sc_hd__xnor2_4 _4449_ (.A(_0456_),
    .B(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__nor2_1 _4450_ (.A(_0455_),
    .B(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__xor2_4 _4451_ (.A(_0455_),
    .B(_0461_),
    .X(_0463_));
 sky130_fd_sc_hd__xor2_4 _4452_ (.A(_0454_),
    .B(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__or2_1 _4453_ (.A(net174),
    .B(net194),
    .X(_0465_));
 sky130_fd_sc_hd__nand2_1 _4454_ (.A(net273),
    .B(net250),
    .Y(_0466_));
 sky130_fd_sc_hd__a2111o_1 _4455_ (.A1(_3381_),
    .A2(_3382_),
    .B1(net250),
    .C1(_3402_),
    .D1(_3365_),
    .X(_0467_));
 sky130_fd_sc_hd__a21o_1 _4456_ (.A1(_0466_),
    .A2(_0467_),
    .B1(_3442_),
    .X(_0468_));
 sky130_fd_sc_hd__or3_1 _4457_ (.A(_3366_),
    .B(_3384_),
    .C(_3400_),
    .X(_0469_));
 sky130_fd_sc_hd__or4_1 _4458_ (.A(_3364_),
    .B(_3383_),
    .C(_3400_),
    .D(net246),
    .X(_0470_));
 sky130_fd_sc_hd__a22oi_1 _4459_ (.A1(net275),
    .A2(net248),
    .B1(_3570_),
    .B2(net274),
    .Y(_0471_));
 sky130_fd_sc_hd__a41o_1 _4460_ (.A1(_0468_),
    .A2(_0469_),
    .A3(_0470_),
    .A4(_0471_),
    .B1(_3406_),
    .X(_0472_));
 sky130_fd_sc_hd__nor2_1 _4461_ (.A(net175),
    .B(net223),
    .Y(_0473_));
 sky130_fd_sc_hd__o22a_1 _4462_ (.A1(net206),
    .A2(net202),
    .B1(net195),
    .B2(net209),
    .X(_0474_));
 sky130_fd_sc_hd__or4_1 _4463_ (.A(net209),
    .B(net206),
    .C(net202),
    .D(net195),
    .X(_0475_));
 sky130_fd_sc_hd__nand2b_1 _4464_ (.A_N(_0474_),
    .B(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__xnor2_1 _4465_ (.A(_0473_),
    .B(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__and2b_1 _4466_ (.A_N(_0465_),
    .B(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__xnor2_2 _4467_ (.A(_0465_),
    .B(_0477_),
    .Y(_0479_));
 sky130_fd_sc_hd__xnor2_2 _4468_ (.A(_0405_),
    .B(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__xor2_4 _4469_ (.A(_0464_),
    .B(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__xnor2_4 _4470_ (.A(_0419_),
    .B(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__xor2_2 _4471_ (.A(_0453_),
    .B(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__a32oi_4 _4472_ (.A1(_0352_),
    .A2(_0362_),
    .A3(_0420_),
    .B1(_0421_),
    .B2(_0385_),
    .Y(_0484_));
 sky130_fd_sc_hd__nand2b_1 _4473_ (.A_N(_0484_),
    .B(_0483_),
    .Y(_0485_));
 sky130_fd_sc_hd__xnor2_2 _4474_ (.A(_0483_),
    .B(_0484_),
    .Y(_0486_));
 sky130_fd_sc_hd__xnor2_2 _4475_ (.A(_0384_),
    .B(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__a21boi_2 _4476_ (.A1(_0336_),
    .A2(_0425_),
    .B1_N(_0424_),
    .Y(_0488_));
 sky130_fd_sc_hd__nor2_1 _4477_ (.A(_0487_),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__xnor2_2 _4478_ (.A(_0487_),
    .B(_0488_),
    .Y(_0490_));
 sky130_fd_sc_hd__xnor2_1 _4479_ (.A(_0427_),
    .B(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__nand3_1 _4480_ (.A(_0429_),
    .B(_0434_),
    .C(_0491_),
    .Y(_0492_));
 sky130_fd_sc_hd__a21o_1 _4481_ (.A1(_0429_),
    .A2(_0434_),
    .B1(_0491_),
    .X(_0493_));
 sky130_fd_sc_hd__and2_1 _4482_ (.A(_0492_),
    .B(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__a21oi_1 _4483_ (.A1(net252),
    .A2(_0435_),
    .B1(_0436_),
    .Y(_0495_));
 sky130_fd_sc_hd__xnor2_1 _4484_ (.A(_0494_),
    .B(_0495_),
    .Y(\mul_wb.reg_p[9] ));
 sky130_fd_sc_hd__a21boi_2 _4485_ (.A1(_0384_),
    .A2(_0486_),
    .B1_N(_0485_),
    .Y(_0496_));
 sky130_fd_sc_hd__a21o_1 _4486_ (.A1(_0381_),
    .A2(_0452_),
    .B1(_0451_),
    .X(_0497_));
 sky130_fd_sc_hd__a21oi_2 _4487_ (.A1(_0454_),
    .A2(_0463_),
    .B1(_0462_),
    .Y(_0498_));
 sky130_fd_sc_hd__a22o_1 _4488_ (.A1(\mul_wb.lob_4.L[12] ),
    .A2(_3495_),
    .B1(_3499_),
    .B2(\mul_wb.lob_4.L[13] ),
    .X(_0499_));
 sky130_fd_sc_hd__and2_1 _4489_ (.A(net244),
    .B(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__nor2_1 _4490_ (.A(_3368_),
    .B(net244),
    .Y(_0501_));
 sky130_fd_sc_hd__a221o_1 _4491_ (.A1(net269),
    .A2(_3543_),
    .B1(_3600_),
    .B2(net271),
    .C1(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__o21ai_1 _4492_ (.A1(_0500_),
    .A2(_0502_),
    .B1(_3488_),
    .Y(_0503_));
 sky130_fd_sc_hd__or2_1 _4493_ (.A(net177),
    .B(net190),
    .X(_0504_));
 sky130_fd_sc_hd__nor2_1 _4494_ (.A(net174),
    .B(net191),
    .Y(_0505_));
 sky130_fd_sc_hd__o22ai_1 _4495_ (.A1(net206),
    .A2(net200),
    .B1(net196),
    .B2(_3683_),
    .Y(_0506_));
 sky130_fd_sc_hd__or4_1 _4496_ (.A(_3683_),
    .B(net206),
    .C(net200),
    .D(net196),
    .X(_0507_));
 sky130_fd_sc_hd__nand2_1 _4497_ (.A(_0506_),
    .B(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__xnor2_2 _4498_ (.A(_0505_),
    .B(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__a21o_1 _4499_ (.A1(_0443_),
    .A2(_0445_),
    .B1(_0446_),
    .X(_0510_));
 sky130_fd_sc_hd__xor2_2 _4500_ (.A(_0509_),
    .B(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__nand2b_1 _4501_ (.A_N(_0504_),
    .B(_0511_),
    .Y(_0512_));
 sky130_fd_sc_hd__xnor2_2 _4502_ (.A(_0504_),
    .B(_0511_),
    .Y(_0513_));
 sky130_fd_sc_hd__nand2b_1 _4503_ (.A_N(_0498_),
    .B(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__xnor2_2 _4504_ (.A(_0498_),
    .B(_0513_),
    .Y(_0515_));
 sky130_fd_sc_hd__nand2b_1 _4505_ (.A_N(_0449_),
    .B(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__xnor2_2 _4506_ (.A(_0449_),
    .B(_0515_),
    .Y(_0517_));
 sky130_fd_sc_hd__o21ai_2 _4507_ (.A1(_0456_),
    .A2(_0460_),
    .B1(_0459_),
    .Y(_0518_));
 sky130_fd_sc_hd__o31a_1 _4508_ (.A1(net175),
    .A2(net223),
    .A3(_0474_),
    .B1(_0475_),
    .X(_0519_));
 sky130_fd_sc_hd__or3b_2 _4509_ (.A(_3527_),
    .B(net198),
    .C_N(_3738_),
    .X(_0520_));
 sky130_fd_sc_hd__nor2_1 _4510_ (.A(net207),
    .B(net195),
    .Y(_0521_));
 sky130_fd_sc_hd__a21oi_2 _4511_ (.A1(net212),
    .A2(net211),
    .B1(net223),
    .Y(_0522_));
 sky130_fd_sc_hd__nand2_1 _4512_ (.A(_0521_),
    .B(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__xnor2_2 _4513_ (.A(_0521_),
    .B(_0522_),
    .Y(_0524_));
 sky130_fd_sc_hd__xnor2_2 _4514_ (.A(_0520_),
    .B(_0524_),
    .Y(_0525_));
 sky130_fd_sc_hd__nor2_1 _4515_ (.A(_0519_),
    .B(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__xor2_2 _4516_ (.A(_0519_),
    .B(_0525_),
    .X(_0527_));
 sky130_fd_sc_hd__xor2_2 _4517_ (.A(_0518_),
    .B(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__or2_1 _4518_ (.A(_3657_),
    .B(net194),
    .X(_0529_));
 sky130_fd_sc_hd__and3_1 _4519_ (.A(net270),
    .B(_3383_),
    .C(_3399_),
    .X(_0530_));
 sky130_fd_sc_hd__a22o_1 _4520_ (.A1(net274),
    .A2(net248),
    .B1(_3444_),
    .B2(net268),
    .X(_0531_));
 sky130_fd_sc_hd__nor2_1 _4521_ (.A(_3367_),
    .B(_3389_),
    .Y(_0532_));
 sky130_fd_sc_hd__and3_1 _4522_ (.A(\mul_wb.lob_4.L[13] ),
    .B(_3389_),
    .C(_3390_),
    .X(_0533_));
 sky130_fd_sc_hd__o21a_1 _4523_ (.A1(_0532_),
    .A2(_0533_),
    .B1(_3396_),
    .X(_0534_));
 sky130_fd_sc_hd__o31ai_4 _4524_ (.A1(_0530_),
    .A2(_0531_),
    .A3(_0534_),
    .B1(net246),
    .Y(_0535_));
 sky130_fd_sc_hd__inv_2 _4525_ (.A(net222),
    .Y(_0536_));
 sky130_fd_sc_hd__or2_1 _4526_ (.A(net175),
    .B(net222),
    .X(_0537_));
 sky130_fd_sc_hd__o22a_1 _4527_ (.A1(net204),
    .A2(net202),
    .B1(net192),
    .B2(net209),
    .X(_0538_));
 sky130_fd_sc_hd__or4_1 _4528_ (.A(net209),
    .B(net204),
    .C(net202),
    .D(net192),
    .X(_0539_));
 sky130_fd_sc_hd__and2b_1 _4529_ (.A_N(_0538_),
    .B(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__xnor2_2 _4530_ (.A(_0537_),
    .B(_0540_),
    .Y(_0541_));
 sky130_fd_sc_hd__and2b_1 _4531_ (.A_N(_0529_),
    .B(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__xnor2_2 _4532_ (.A(_0529_),
    .B(_0541_),
    .Y(_0543_));
 sky130_fd_sc_hd__and2_1 _4533_ (.A(_0478_),
    .B(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__xor2_2 _4534_ (.A(_0478_),
    .B(_0543_),
    .X(_0545_));
 sky130_fd_sc_hd__xnor2_2 _4535_ (.A(_0528_),
    .B(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__a32o_1 _4536_ (.A1(_0392_),
    .A2(_0404_),
    .A3(_0479_),
    .B1(_0480_),
    .B2(_0464_),
    .X(_0547_));
 sky130_fd_sc_hd__nand2b_1 _4537_ (.A_N(_0546_),
    .B(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__xnor2_2 _4538_ (.A(_0546_),
    .B(_0547_),
    .Y(_0549_));
 sky130_fd_sc_hd__xor2_2 _4539_ (.A(_0517_),
    .B(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__a32oi_4 _4540_ (.A1(_0407_),
    .A2(_0418_),
    .A3(_0481_),
    .B1(_0482_),
    .B2(_0453_),
    .Y(_0551_));
 sky130_fd_sc_hd__and2b_1 _4541_ (.A_N(_0551_),
    .B(_0550_),
    .X(_0552_));
 sky130_fd_sc_hd__xnor2_2 _4542_ (.A(_0550_),
    .B(_0551_),
    .Y(_0553_));
 sky130_fd_sc_hd__xor2_2 _4543_ (.A(_0497_),
    .B(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__nand2b_1 _4544_ (.A_N(_0496_),
    .B(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__xnor2_2 _4545_ (.A(_0496_),
    .B(_0554_),
    .Y(_0556_));
 sky130_fd_sc_hd__nand2_1 _4546_ (.A(_0489_),
    .B(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__xnor2_2 _4547_ (.A(_0489_),
    .B(_0556_),
    .Y(_0558_));
 sky130_fd_sc_hd__a211o_1 _4548_ (.A1(_0373_),
    .A2(_0432_),
    .B1(_0491_),
    .C1(_0430_),
    .X(_0559_));
 sky130_fd_sc_hd__a21o_1 _4549_ (.A1(_0427_),
    .A2(_0429_),
    .B1(_0490_),
    .X(_0560_));
 sky130_fd_sc_hd__a21o_1 _4550_ (.A1(_0559_),
    .A2(_0560_),
    .B1(_0558_),
    .X(_0561_));
 sky130_fd_sc_hd__nand3_1 _4551_ (.A(_0558_),
    .B(_0559_),
    .C(_0560_),
    .Y(_0562_));
 sky130_fd_sc_hd__and2_2 _4552_ (.A(_0561_),
    .B(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__a2111o_2 _4553_ (.A1(_0492_),
    .A2(_0493_),
    .B1(_0322_),
    .C1(_0375_),
    .D1(_0435_),
    .X(_0564_));
 sky130_fd_sc_hd__nand2_1 _4554_ (.A(net252),
    .B(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__xnor2_1 _4555_ (.A(_0563_),
    .B(_0565_),
    .Y(\mul_wb.reg_p[10] ));
 sky130_fd_sc_hd__or2_1 _4556_ (.A(_0563_),
    .B(_0564_),
    .X(_0566_));
 sky130_fd_sc_hd__nand2_1 _4557_ (.A(net252),
    .B(_0566_),
    .Y(_0567_));
 sky130_fd_sc_hd__nand2_1 _4558_ (.A(_0514_),
    .B(_0516_),
    .Y(_0568_));
 sky130_fd_sc_hd__a21bo_1 _4559_ (.A1(_0509_),
    .A2(_0510_),
    .B1_N(_0512_),
    .X(_0569_));
 sky130_fd_sc_hd__a21oi_2 _4560_ (.A1(_0518_),
    .A2(_0527_),
    .B1(_0526_),
    .Y(_0570_));
 sky130_fd_sc_hd__nor2_1 _4561_ (.A(net174),
    .B(net190),
    .Y(_0571_));
 sky130_fd_sc_hd__or2_1 _4562_ (.A(_3657_),
    .B(net191),
    .X(_0572_));
 sky130_fd_sc_hd__o22ai_1 _4563_ (.A1(net204),
    .A2(net200),
    .B1(net196),
    .B2(net206),
    .Y(_0573_));
 sky130_fd_sc_hd__or4_1 _4564_ (.A(net206),
    .B(net204),
    .C(net200),
    .D(net196),
    .X(_0574_));
 sky130_fd_sc_hd__nand2_1 _4565_ (.A(_0573_),
    .B(_0574_),
    .Y(_0575_));
 sky130_fd_sc_hd__xnor2_2 _4566_ (.A(_0572_),
    .B(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__o31a_1 _4567_ (.A1(net174),
    .A2(net191),
    .A3(_0508_),
    .B1(_0507_),
    .X(_0577_));
 sky130_fd_sc_hd__nor2_1 _4568_ (.A(_0576_),
    .B(_0577_),
    .Y(_0578_));
 sky130_fd_sc_hd__xor2_2 _4569_ (.A(_0576_),
    .B(_0577_),
    .X(_0579_));
 sky130_fd_sc_hd__xor2_2 _4570_ (.A(_0571_),
    .B(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__nand2b_1 _4571_ (.A_N(_0570_),
    .B(_0580_),
    .Y(_0581_));
 sky130_fd_sc_hd__xnor2_2 _4572_ (.A(_0570_),
    .B(_0580_),
    .Y(_0582_));
 sky130_fd_sc_hd__xor2_2 _4573_ (.A(_0569_),
    .B(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__o21ai_2 _4574_ (.A1(_0520_),
    .A2(_0524_),
    .B1(_0523_),
    .Y(_0584_));
 sky130_fd_sc_hd__o21a_1 _4575_ (.A1(_0537_),
    .A2(_0538_),
    .B1(_0539_),
    .X(_0585_));
 sky130_fd_sc_hd__or3b_2 _4576_ (.A(_3527_),
    .B(net195),
    .C_N(_3738_),
    .X(_0586_));
 sky130_fd_sc_hd__nor2_1 _4577_ (.A(net207),
    .B(net192),
    .Y(_0587_));
 sky130_fd_sc_hd__a21oi_2 _4578_ (.A1(net212),
    .A2(net211),
    .B1(net222),
    .Y(_0588_));
 sky130_fd_sc_hd__nand2_1 _4579_ (.A(_0587_),
    .B(_0588_),
    .Y(_0589_));
 sky130_fd_sc_hd__xnor2_2 _4580_ (.A(_0587_),
    .B(_0588_),
    .Y(_0590_));
 sky130_fd_sc_hd__xnor2_2 _4581_ (.A(_0586_),
    .B(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__nor2_1 _4582_ (.A(_0585_),
    .B(_0591_),
    .Y(_0592_));
 sky130_fd_sc_hd__xor2_2 _4583_ (.A(_0585_),
    .B(_0591_),
    .X(_0593_));
 sky130_fd_sc_hd__xor2_2 _4584_ (.A(_0584_),
    .B(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__a22o_1 _4585_ (.A1(net273),
    .A2(net248),
    .B1(_3568_),
    .B2(net270),
    .X(_0595_));
 sky130_fd_sc_hd__a22o_1 _4586_ (.A1(net268),
    .A2(_3399_),
    .B1(_3570_),
    .B2(net272),
    .X(_0596_));
 sky130_fd_sc_hd__o21a_1 _4587_ (.A1(_0595_),
    .A2(_0596_),
    .B1(_3383_),
    .X(_0597_));
 sky130_fd_sc_hd__o21ai_4 _4588_ (.A1(_0595_),
    .A2(_0596_),
    .B1(_3383_),
    .Y(_0598_));
 sky130_fd_sc_hd__nor2_1 _4589_ (.A(net175),
    .B(net221),
    .Y(_0599_));
 sky130_fd_sc_hd__o22a_1 _4590_ (.A1(net202),
    .A2(net198),
    .B1(net223),
    .B2(net209),
    .X(_0600_));
 sky130_fd_sc_hd__or4_1 _4591_ (.A(net209),
    .B(net202),
    .C(net198),
    .D(net223),
    .X(_0601_));
 sky130_fd_sc_hd__nand2b_1 _4592_ (.A_N(_0600_),
    .B(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__xnor2_2 _4593_ (.A(_0599_),
    .B(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__a22o_1 _4594_ (.A1(\mul_wb.lob_4.L[13] ),
    .A2(_3589_),
    .B1(_3601_),
    .B2(net270),
    .X(_0604_));
 sky130_fd_sc_hd__a32o_1 _4595_ (.A1(net268),
    .A2(_3497_),
    .A3(_3513_),
    .B1(\mul_wb.lob_4.L[12] ),
    .B2(net245),
    .X(_0605_));
 sky130_fd_sc_hd__o21a_1 _4596_ (.A1(_0604_),
    .A2(_0605_),
    .B1(_3487_),
    .X(_0606_));
 sky130_fd_sc_hd__o21ai_2 _4597_ (.A1(_0604_),
    .A2(_0605_),
    .B1(_3487_),
    .Y(_0607_));
 sky130_fd_sc_hd__nor2_1 _4598_ (.A(net177),
    .B(net220),
    .Y(_0608_));
 sky130_fd_sc_hd__nor2_1 _4599_ (.A(net208),
    .B(net194),
    .Y(_0609_));
 sky130_fd_sc_hd__or3b_1 _4600_ (.A(_3475_),
    .B(net220),
    .C_N(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__xor2_2 _4601_ (.A(_0608_),
    .B(_0609_),
    .X(_0611_));
 sky130_fd_sc_hd__nand2_1 _4602_ (.A(_0603_),
    .B(_0611_),
    .Y(_0612_));
 sky130_fd_sc_hd__xor2_2 _4603_ (.A(_0603_),
    .B(_0611_),
    .X(_0613_));
 sky130_fd_sc_hd__and2_1 _4604_ (.A(_0542_),
    .B(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__xor2_2 _4605_ (.A(_0542_),
    .B(_0613_),
    .X(_0615_));
 sky130_fd_sc_hd__xnor2_2 _4606_ (.A(_0594_),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__a21oi_2 _4607_ (.A1(_0528_),
    .A2(_0545_),
    .B1(_0544_),
    .Y(_0617_));
 sky130_fd_sc_hd__nor2_1 _4608_ (.A(_0616_),
    .B(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__xor2_2 _4609_ (.A(_0616_),
    .B(_0617_),
    .X(_0619_));
 sky130_fd_sc_hd__xnor2_2 _4610_ (.A(_0583_),
    .B(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__a21boi_2 _4611_ (.A1(_0517_),
    .A2(_0549_),
    .B1_N(_0548_),
    .Y(_0621_));
 sky130_fd_sc_hd__nor2_1 _4612_ (.A(_0620_),
    .B(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__xor2_2 _4613_ (.A(_0620_),
    .B(_0621_),
    .X(_0623_));
 sky130_fd_sc_hd__xnor2_2 _4614_ (.A(_0568_),
    .B(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__a21oi_2 _4615_ (.A1(_0497_),
    .A2(_0553_),
    .B1(_0552_),
    .Y(_0625_));
 sky130_fd_sc_hd__nor2_1 _4616_ (.A(_0624_),
    .B(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__xnor2_2 _4617_ (.A(_0624_),
    .B(_0625_),
    .Y(_0627_));
 sky130_fd_sc_hd__xnor2_2 _4618_ (.A(_0555_),
    .B(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__nand3_2 _4619_ (.A(_0557_),
    .B(_0561_),
    .C(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__a21o_1 _4620_ (.A1(_0557_),
    .A2(_0561_),
    .B1(_0628_),
    .X(_0630_));
 sky130_fd_sc_hd__and2_1 _4621_ (.A(_0629_),
    .B(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__xnor2_1 _4622_ (.A(_0567_),
    .B(_0631_),
    .Y(\mul_wb.reg_p[11] ));
 sky130_fd_sc_hd__a21o_1 _4623_ (.A1(_0568_),
    .A2(_0623_),
    .B1(_0622_),
    .X(_0632_));
 sky130_fd_sc_hd__a21bo_1 _4624_ (.A1(_0569_),
    .A2(_0582_),
    .B1_N(_0581_),
    .X(_0633_));
 sky130_fd_sc_hd__a21o_1 _4625_ (.A1(_0571_),
    .A2(_0579_),
    .B1(_0578_),
    .X(_0634_));
 sky130_fd_sc_hd__a21o_1 _4626_ (.A1(_0584_),
    .A2(_0593_),
    .B1(_0592_),
    .X(_0635_));
 sky130_fd_sc_hd__o21ai_1 _4627_ (.A1(net272),
    .A2(_3484_),
    .B1(net243),
    .Y(_0636_));
 sky130_fd_sc_hd__a221o_2 _4628_ (.A1(_3364_),
    .A2(_3542_),
    .B1(_3589_),
    .B2(_3365_),
    .C1(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__or4_2 _4629_ (.A(_3475_),
    .B(_3657_),
    .C(net190),
    .D(net219),
    .X(_0638_));
 sky130_fd_sc_hd__o22ai_2 _4630_ (.A1(_3657_),
    .A2(net190),
    .B1(net219),
    .B2(_3475_),
    .Y(_0639_));
 sky130_fd_sc_hd__nand2_1 _4631_ (.A(_0638_),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__or2_1 _4632_ (.A(_3683_),
    .B(net191),
    .X(_0641_));
 sky130_fd_sc_hd__o22a_1 _4633_ (.A1(net200),
    .A2(net198),
    .B1(net196),
    .B2(net204),
    .X(_0642_));
 sky130_fd_sc_hd__or4_1 _4634_ (.A(net204),
    .B(net200),
    .C(net198),
    .D(net196),
    .X(_0643_));
 sky130_fd_sc_hd__and2b_1 _4635_ (.A_N(_0642_),
    .B(_0643_),
    .X(_0644_));
 sky130_fd_sc_hd__xnor2_1 _4636_ (.A(_0641_),
    .B(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__o21a_1 _4637_ (.A1(_0572_),
    .A2(_0575_),
    .B1(_0574_),
    .X(_0646_));
 sky130_fd_sc_hd__and2b_1 _4638_ (.A_N(_0646_),
    .B(_0645_),
    .X(_0647_));
 sky130_fd_sc_hd__xnor2_1 _4639_ (.A(_0645_),
    .B(_0646_),
    .Y(_0648_));
 sky130_fd_sc_hd__xnor2_1 _4640_ (.A(_0640_),
    .B(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__xnor2_1 _4641_ (.A(_0635_),
    .B(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__and2b_1 _4642_ (.A_N(_0650_),
    .B(_0634_),
    .X(_0651_));
 sky130_fd_sc_hd__xnor2_1 _4643_ (.A(_0634_),
    .B(_0650_),
    .Y(_0652_));
 sky130_fd_sc_hd__o21ai_1 _4644_ (.A1(_0586_),
    .A2(_0590_),
    .B1(_0589_),
    .Y(_0653_));
 sky130_fd_sc_hd__o31a_1 _4645_ (.A1(net175),
    .A2(net221),
    .A3(_0600_),
    .B1(_0601_),
    .X(_0654_));
 sky130_fd_sc_hd__nor2_1 _4646_ (.A(net207),
    .B(net223),
    .Y(_0655_));
 sky130_fd_sc_hd__a21oi_2 _4647_ (.A1(net212),
    .A2(net211),
    .B1(net221),
    .Y(_0656_));
 sky130_fd_sc_hd__nand2_1 _4648_ (.A(_0655_),
    .B(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__xnor2_2 _4649_ (.A(_0655_),
    .B(_0656_),
    .Y(_0658_));
 sky130_fd_sc_hd__or3b_2 _4650_ (.A(_3527_),
    .B(net192),
    .C_N(_3738_),
    .X(_0659_));
 sky130_fd_sc_hd__xnor2_2 _4651_ (.A(_0658_),
    .B(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__nor2_1 _4652_ (.A(_0654_),
    .B(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__nand2_1 _4653_ (.A(_0654_),
    .B(_0660_),
    .Y(_0662_));
 sky130_fd_sc_hd__xnor2_1 _4654_ (.A(_0654_),
    .B(_0660_),
    .Y(_0663_));
 sky130_fd_sc_hd__xnor2_1 _4655_ (.A(_0653_),
    .B(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__or3_1 _4656_ (.A(net270),
    .B(_3389_),
    .C(net248),
    .X(_0665_));
 sky130_fd_sc_hd__o21a_1 _4657_ (.A1(net272),
    .A2(_3396_),
    .B1(net250),
    .X(_0666_));
 sky130_fd_sc_hd__o211ai_4 _4658_ (.A1(net268),
    .A2(_3442_),
    .B1(_0665_),
    .C1(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__inv_2 _4659_ (.A(net227),
    .Y(_0668_));
 sky130_fd_sc_hd__nor2_1 _4660_ (.A(net175),
    .B(net227),
    .Y(_0669_));
 sky130_fd_sc_hd__o22ai_1 _4661_ (.A1(net202),
    .A2(net195),
    .B1(net222),
    .B2(net210),
    .Y(_0670_));
 sky130_fd_sc_hd__or4_1 _4662_ (.A(net210),
    .B(net202),
    .C(net195),
    .D(net222),
    .X(_0671_));
 sky130_fd_sc_hd__nand2_1 _4663_ (.A(_0670_),
    .B(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__xnor2_1 _4664_ (.A(_0669_),
    .B(_0672_),
    .Y(_0673_));
 sky130_fd_sc_hd__a21o_1 _4665_ (.A1(_3583_),
    .A2(_3586_),
    .B1(net220),
    .X(_0674_));
 sky130_fd_sc_hd__nor2_1 _4666_ (.A(net206),
    .B(net194),
    .Y(_0675_));
 sky130_fd_sc_hd__or3_1 _4667_ (.A(net206),
    .B(net194),
    .C(_0674_),
    .X(_0676_));
 sky130_fd_sc_hd__xnor2_1 _4668_ (.A(_0674_),
    .B(_0675_),
    .Y(_0677_));
 sky130_fd_sc_hd__xnor2_1 _4669_ (.A(_0610_),
    .B(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__xnor2_1 _4670_ (.A(_0673_),
    .B(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__nor2_1 _4671_ (.A(_0612_),
    .B(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__xor2_1 _4672_ (.A(_0612_),
    .B(_0679_),
    .X(_0681_));
 sky130_fd_sc_hd__xnor2_1 _4673_ (.A(_0664_),
    .B(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__a21o_1 _4674_ (.A1(_0594_),
    .A2(_0615_),
    .B1(_0614_),
    .X(_0683_));
 sky130_fd_sc_hd__and2b_1 _4675_ (.A_N(_0682_),
    .B(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__xnor2_1 _4676_ (.A(_0682_),
    .B(_0683_),
    .Y(_0685_));
 sky130_fd_sc_hd__xnor2_1 _4677_ (.A(_0652_),
    .B(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__a21oi_1 _4678_ (.A1(_0583_),
    .A2(_0619_),
    .B1(_0618_),
    .Y(_0687_));
 sky130_fd_sc_hd__xnor2_1 _4679_ (.A(_0686_),
    .B(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__nand2b_1 _4680_ (.A_N(_0688_),
    .B(_0633_),
    .Y(_0689_));
 sky130_fd_sc_hd__xor2_1 _4681_ (.A(_0633_),
    .B(_0688_),
    .X(_0690_));
 sky130_fd_sc_hd__nand2b_2 _4682_ (.A_N(_0690_),
    .B(_0632_),
    .Y(_0691_));
 sky130_fd_sc_hd__xnor2_1 _4683_ (.A(_0632_),
    .B(_0690_),
    .Y(_0692_));
 sky130_fd_sc_hd__nand2_1 _4684_ (.A(_0626_),
    .B(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hd__or2_1 _4685_ (.A(_0626_),
    .B(_0692_),
    .X(_0694_));
 sky130_fd_sc_hd__and2_2 _4686_ (.A(_0693_),
    .B(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__inv_2 _4687_ (.A(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__a21o_1 _4688_ (.A1(_0555_),
    .A2(_0557_),
    .B1(_0627_),
    .X(_0697_));
 sky130_fd_sc_hd__a2111o_1 _4689_ (.A1(_0427_),
    .A2(_0429_),
    .B1(_0490_),
    .C1(_0558_),
    .D1(_0628_),
    .X(_0698_));
 sky130_fd_sc_hd__o311a_4 _4690_ (.A1(_0558_),
    .A2(_0559_),
    .A3(_0628_),
    .B1(_0697_),
    .C1(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__xnor2_4 _4691_ (.A(_0695_),
    .B(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__o21a_1 _4692_ (.A1(_0566_),
    .A2(_0631_),
    .B1(net252),
    .X(_0701_));
 sky130_fd_sc_hd__xor2_1 _4693_ (.A(_0700_),
    .B(_0701_),
    .X(\mul_wb.reg_p[12] ));
 sky130_fd_sc_hd__a2111oi_4 _4694_ (.A1(_0629_),
    .A2(_0630_),
    .B1(_0700_),
    .C1(_0564_),
    .D1(_0563_),
    .Y(_0702_));
 sky130_fd_sc_hd__or2_1 _4695_ (.A(_3620_),
    .B(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__o21ai_2 _4696_ (.A1(_0696_),
    .A2(_0699_),
    .B1(_0693_),
    .Y(_0704_));
 sky130_fd_sc_hd__a21oi_1 _4697_ (.A1(_0635_),
    .A2(_0649_),
    .B1(_0651_),
    .Y(_0705_));
 sky130_fd_sc_hd__or2_1 _4698_ (.A(_0638_),
    .B(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__nand2_1 _4699_ (.A(_0638_),
    .B(_0705_),
    .Y(_0707_));
 sky130_fd_sc_hd__and2_1 _4700_ (.A(_0706_),
    .B(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__a31oi_2 _4701_ (.A1(_0638_),
    .A2(_0639_),
    .A3(_0648_),
    .B1(_0647_),
    .Y(_0709_));
 sky130_fd_sc_hd__a21o_1 _4702_ (.A1(_0653_),
    .A2(_0662_),
    .B1(_0661_),
    .X(_0710_));
 sky130_fd_sc_hd__o22a_1 _4703_ (.A1(_3683_),
    .A2(net190),
    .B1(net219),
    .B2(net174),
    .X(_0711_));
 sky130_fd_sc_hd__or4_1 _4704_ (.A(_3587_),
    .B(_3683_),
    .C(net190),
    .D(net219),
    .X(_0712_));
 sky130_fd_sc_hd__and2b_1 _4705_ (.A_N(_0711_),
    .B(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__a22o_1 _4706_ (.A1(net271),
    .A2(net245),
    .B1(_3513_),
    .B2(net268),
    .X(_0714_));
 sky130_fd_sc_hd__nand2_2 _4707_ (.A(_3495_),
    .B(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__nor2_1 _4708_ (.A(_3475_),
    .B(net217),
    .Y(_0716_));
 sky130_fd_sc_hd__xnor2_2 _4709_ (.A(_0713_),
    .B(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__o22ai_1 _4710_ (.A1(net198),
    .A2(net196),
    .B1(net195),
    .B2(net200),
    .Y(_0718_));
 sky130_fd_sc_hd__or4_1 _4711_ (.A(net200),
    .B(net198),
    .C(net196),
    .D(net195),
    .X(_0719_));
 sky130_fd_sc_hd__nand2_1 _4712_ (.A(_0718_),
    .B(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__or2_1 _4713_ (.A(net206),
    .B(net191),
    .X(_0721_));
 sky130_fd_sc_hd__xnor2_2 _4714_ (.A(_0720_),
    .B(_0721_),
    .Y(_0722_));
 sky130_fd_sc_hd__o21a_1 _4715_ (.A1(_0641_),
    .A2(_0642_),
    .B1(_0643_),
    .X(_0723_));
 sky130_fd_sc_hd__or2_1 _4716_ (.A(_0722_),
    .B(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__xnor2_2 _4717_ (.A(_0722_),
    .B(_0723_),
    .Y(_0725_));
 sky130_fd_sc_hd__xor2_1 _4718_ (.A(_0717_),
    .B(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__and2_1 _4719_ (.A(_0710_),
    .B(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__xor2_1 _4720_ (.A(_0710_),
    .B(_0726_),
    .X(_0728_));
 sky130_fd_sc_hd__and2b_1 _4721_ (.A_N(_0709_),
    .B(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__xnor2_1 _4722_ (.A(_0709_),
    .B(_0728_),
    .Y(_0730_));
 sky130_fd_sc_hd__o21ai_1 _4723_ (.A1(_0658_),
    .A2(_0659_),
    .B1(_0657_),
    .Y(_0731_));
 sky130_fd_sc_hd__o31a_1 _4724_ (.A1(net175),
    .A2(_0667_),
    .A3(_0672_),
    .B1(_0671_),
    .X(_0732_));
 sky130_fd_sc_hd__nor2_1 _4725_ (.A(net207),
    .B(net222),
    .Y(_0733_));
 sky130_fd_sc_hd__a21oi_2 _4726_ (.A1(net212),
    .A2(net211),
    .B1(_0667_),
    .Y(_0734_));
 sky130_fd_sc_hd__nand2_1 _4727_ (.A(_0733_),
    .B(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__xnor2_2 _4728_ (.A(_0733_),
    .B(_0734_),
    .Y(_0736_));
 sky130_fd_sc_hd__or3b_2 _4729_ (.A(_3527_),
    .B(net223),
    .C_N(_3738_),
    .X(_0737_));
 sky130_fd_sc_hd__xnor2_1 _4730_ (.A(_0736_),
    .B(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__nor2_1 _4731_ (.A(_0732_),
    .B(_0738_),
    .Y(_0739_));
 sky130_fd_sc_hd__xor2_1 _4732_ (.A(_0732_),
    .B(_0738_),
    .X(_0740_));
 sky130_fd_sc_hd__xnor2_1 _4733_ (.A(_0731_),
    .B(_0740_),
    .Y(_0741_));
 sky130_fd_sc_hd__a21oi_1 _4734_ (.A1(_3648_),
    .A2(_3656_),
    .B1(net220),
    .Y(_0742_));
 sky130_fd_sc_hd__or2_1 _4735_ (.A(net204),
    .B(net194),
    .X(_0743_));
 sky130_fd_sc_hd__or3_2 _4736_ (.A(_3657_),
    .B(net220),
    .C(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__xnor2_1 _4737_ (.A(_0742_),
    .B(_0743_),
    .Y(_0745_));
 sky130_fd_sc_hd__nand2b_1 _4738_ (.A_N(_0676_),
    .B(_0745_),
    .Y(_0746_));
 sky130_fd_sc_hd__xnor2_1 _4739_ (.A(_0676_),
    .B(_0745_),
    .Y(_0747_));
 sky130_fd_sc_hd__o22ai_1 _4740_ (.A1(net203),
    .A2(net192),
    .B1(net221),
    .B2(net210),
    .Y(_0748_));
 sky130_fd_sc_hd__or4_1 _4741_ (.A(net209),
    .B(net203),
    .C(net192),
    .D(net221),
    .X(_0749_));
 sky130_fd_sc_hd__nand2_1 _4742_ (.A(_0748_),
    .B(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__a22o_1 _4743_ (.A1(net270),
    .A2(net249),
    .B1(_3398_),
    .B2(net268),
    .X(_0751_));
 sky130_fd_sc_hd__and2_2 _4744_ (.A(_3388_),
    .B(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__nand2_2 _4745_ (.A(_3388_),
    .B(_0751_),
    .Y(_0753_));
 sky130_fd_sc_hd__nor2_1 _4746_ (.A(net175),
    .B(net216),
    .Y(_0754_));
 sky130_fd_sc_hd__or3_1 _4747_ (.A(net176),
    .B(_0750_),
    .C(net216),
    .X(_0755_));
 sky130_fd_sc_hd__xnor2_1 _4748_ (.A(_0750_),
    .B(_0754_),
    .Y(_0756_));
 sky130_fd_sc_hd__xnor2_1 _4749_ (.A(_0747_),
    .B(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__a32o_1 _4750_ (.A1(_0608_),
    .A2(_0609_),
    .A3(_0677_),
    .B1(_0678_),
    .B2(_0673_),
    .X(_0758_));
 sky130_fd_sc_hd__and2b_1 _4751_ (.A_N(_0757_),
    .B(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__xor2_1 _4752_ (.A(_0757_),
    .B(_0758_),
    .X(_0760_));
 sky130_fd_sc_hd__xnor2_1 _4753_ (.A(_0741_),
    .B(_0760_),
    .Y(_0761_));
 sky130_fd_sc_hd__a21oi_1 _4754_ (.A1(_0664_),
    .A2(_0681_),
    .B1(_0680_),
    .Y(_0762_));
 sky130_fd_sc_hd__nor2_1 _4755_ (.A(_0761_),
    .B(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__xor2_1 _4756_ (.A(_0761_),
    .B(_0762_),
    .X(_0764_));
 sky130_fd_sc_hd__xnor2_1 _4757_ (.A(_0730_),
    .B(_0764_),
    .Y(_0765_));
 sky130_fd_sc_hd__a21oi_1 _4758_ (.A1(_0652_),
    .A2(_0685_),
    .B1(_0684_),
    .Y(_0766_));
 sky130_fd_sc_hd__nor2_1 _4759_ (.A(_0765_),
    .B(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__nand2_1 _4760_ (.A(_0765_),
    .B(_0766_),
    .Y(_0768_));
 sky130_fd_sc_hd__and2b_1 _4761_ (.A_N(_0767_),
    .B(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__xnor2_1 _4762_ (.A(_0708_),
    .B(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__o21a_1 _4763_ (.A1(_0686_),
    .A2(_0687_),
    .B1(_0689_),
    .X(_0771_));
 sky130_fd_sc_hd__nor2_1 _4764_ (.A(_0770_),
    .B(_0771_),
    .Y(_0772_));
 sky130_fd_sc_hd__and2_1 _4765_ (.A(_0770_),
    .B(_0771_),
    .X(_0773_));
 sky130_fd_sc_hd__or2_2 _4766_ (.A(_0772_),
    .B(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__xnor2_4 _4767_ (.A(_0691_),
    .B(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__xnor2_4 _4768_ (.A(_0704_),
    .B(_0775_),
    .Y(_0776_));
 sky130_fd_sc_hd__xnor2_2 _4769_ (.A(_0703_),
    .B(_0776_),
    .Y(\mul_wb.reg_p[13] ));
 sky130_fd_sc_hd__a21boi_1 _4770_ (.A1(_0713_),
    .A2(_0716_),
    .B1_N(_0712_),
    .Y(_0777_));
 sky130_fd_sc_hd__o21ba_1 _4771_ (.A1(_0727_),
    .A2(_0729_),
    .B1_N(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__or3b_1 _4772_ (.A(_0727_),
    .B(_0729_),
    .C_N(_0777_),
    .X(_0779_));
 sky130_fd_sc_hd__and2b_1 _4773_ (.A_N(_0778_),
    .B(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__o21ai_4 _4774_ (.A1(_0717_),
    .A2(_0725_),
    .B1(_0724_),
    .Y(_0781_));
 sky130_fd_sc_hd__a21o_2 _4775_ (.A1(_0731_),
    .A2(_0740_),
    .B1(_0739_),
    .X(_0782_));
 sky130_fd_sc_hd__o22ai_2 _4776_ (.A1(_3722_),
    .A2(net190),
    .B1(net219),
    .B2(net173),
    .Y(_0783_));
 sky130_fd_sc_hd__or4_1 _4777_ (.A(net173),
    .B(_3722_),
    .C(net190),
    .D(net219),
    .X(_0784_));
 sky130_fd_sc_hd__nand2_2 _4778_ (.A(_0783_),
    .B(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__nor2_2 _4779_ (.A(_3587_),
    .B(net217),
    .Y(_0786_));
 sky130_fd_sc_hd__xor2_4 _4780_ (.A(_0785_),
    .B(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__o22a_1 _4781_ (.A1(net197),
    .A2(net195),
    .B1(net192),
    .B2(net201),
    .X(_0788_));
 sky130_fd_sc_hd__or4_1 _4782_ (.A(net201),
    .B(net196),
    .C(net195),
    .D(net192),
    .X(_0789_));
 sky130_fd_sc_hd__and2b_1 _4783_ (.A_N(_0788_),
    .B(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__nor2_2 _4784_ (.A(net204),
    .B(net191),
    .Y(_0791_));
 sky130_fd_sc_hd__xnor2_4 _4785_ (.A(_0790_),
    .B(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__o21a_2 _4786_ (.A1(_0720_),
    .A2(_0721_),
    .B1(_0719_),
    .X(_0793_));
 sky130_fd_sc_hd__xor2_4 _4787_ (.A(_0792_),
    .B(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__nand2b_1 _4788_ (.A_N(_0787_),
    .B(_0794_),
    .Y(_0795_));
 sky130_fd_sc_hd__xnor2_4 _4789_ (.A(_0787_),
    .B(_0794_),
    .Y(_0796_));
 sky130_fd_sc_hd__and2_1 _4790_ (.A(_0782_),
    .B(_0796_),
    .X(_0797_));
 sky130_fd_sc_hd__xnor2_4 _4791_ (.A(_0782_),
    .B(_0796_),
    .Y(_0798_));
 sky130_fd_sc_hd__and2b_1 _4792_ (.A_N(_0798_),
    .B(_0781_),
    .X(_0799_));
 sky130_fd_sc_hd__xnor2_4 _4793_ (.A(_0781_),
    .B(_0798_),
    .Y(_0800_));
 sky130_fd_sc_hd__o21ai_4 _4794_ (.A1(_0736_),
    .A2(_0737_),
    .B1(_0735_),
    .Y(_0801_));
 sky130_fd_sc_hd__inv_2 _4795_ (.A(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__or2_1 _4796_ (.A(net207),
    .B(net221),
    .X(_0803_));
 sky130_fd_sc_hd__a21oi_1 _4797_ (.A1(net212),
    .A2(net211),
    .B1(net216),
    .Y(_0804_));
 sky130_fd_sc_hd__or3_1 _4798_ (.A(_3614_),
    .B(_0753_),
    .C(_0803_),
    .X(_0805_));
 sky130_fd_sc_hd__xnor2_1 _4799_ (.A(_0803_),
    .B(_0804_),
    .Y(_0806_));
 sky130_fd_sc_hd__and3_1 _4800_ (.A(_3526_),
    .B(_3738_),
    .C(_0536_),
    .X(_0807_));
 sky130_fd_sc_hd__xnor2_1 _4801_ (.A(_0806_),
    .B(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__a21oi_1 _4802_ (.A1(_0749_),
    .A2(_0755_),
    .B1(_0808_),
    .Y(_0809_));
 sky130_fd_sc_hd__and3_1 _4803_ (.A(_0749_),
    .B(_0755_),
    .C(_0808_),
    .X(_0810_));
 sky130_fd_sc_hd__or2_2 _4804_ (.A(_0809_),
    .B(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__xnor2_4 _4805_ (.A(_0801_),
    .B(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__or2_2 _4806_ (.A(net203),
    .B(net223),
    .X(_0813_));
 sky130_fd_sc_hd__or2_2 _4807_ (.A(net210),
    .B(_0667_),
    .X(_0814_));
 sky130_fd_sc_hd__xnor2_4 _4808_ (.A(_0813_),
    .B(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__nand2_2 _4809_ (.A(net268),
    .B(net249),
    .Y(_0816_));
 sky130_fd_sc_hd__or2_2 _4810_ (.A(net175),
    .B(net237),
    .X(_0817_));
 sky130_fd_sc_hd__xnor2_4 _4811_ (.A(_0815_),
    .B(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__nor2_2 _4812_ (.A(net198),
    .B(net194),
    .Y(_0819_));
 sky130_fd_sc_hd__or2_2 _4813_ (.A(net208),
    .B(net220),
    .X(_0820_));
 sky130_fd_sc_hd__nor2_2 _4814_ (.A(_3364_),
    .B(net244),
    .Y(_0821_));
 sky130_fd_sc_hd__nand2_8 _4815_ (.A(net269),
    .B(net245),
    .Y(_0822_));
 sky130_fd_sc_hd__a31oi_4 _4816_ (.A1(_3455_),
    .A2(_3467_),
    .A3(_3474_),
    .B1(_0822_),
    .Y(_0823_));
 sky130_fd_sc_hd__and2b_1 _4817_ (.A_N(_0820_),
    .B(_0823_),
    .X(_0824_));
 sky130_fd_sc_hd__xnor2_4 _4818_ (.A(_0820_),
    .B(_0823_),
    .Y(_0825_));
 sky130_fd_sc_hd__xnor2_4 _4819_ (.A(_0819_),
    .B(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__nor2_1 _4820_ (.A(_0744_),
    .B(_0826_),
    .Y(_0827_));
 sky130_fd_sc_hd__xnor2_4 _4821_ (.A(_0744_),
    .B(_0826_),
    .Y(_0828_));
 sky130_fd_sc_hd__xnor2_4 _4822_ (.A(_0818_),
    .B(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__a21bo_2 _4823_ (.A1(_0747_),
    .A2(_0756_),
    .B1_N(_0746_),
    .X(_0830_));
 sky130_fd_sc_hd__nand2b_1 _4824_ (.A_N(_0829_),
    .B(_0830_),
    .Y(_0831_));
 sky130_fd_sc_hd__xnor2_4 _4825_ (.A(_0829_),
    .B(_0830_),
    .Y(_0832_));
 sky130_fd_sc_hd__xor2_4 _4826_ (.A(_0812_),
    .B(_0832_),
    .X(_0833_));
 sky130_fd_sc_hd__o21ba_2 _4827_ (.A1(_0741_),
    .A2(_0760_),
    .B1_N(_0759_),
    .X(_0834_));
 sky130_fd_sc_hd__and2b_1 _4828_ (.A_N(_0834_),
    .B(_0833_),
    .X(_0835_));
 sky130_fd_sc_hd__xnor2_4 _4829_ (.A(_0833_),
    .B(_0834_),
    .Y(_0836_));
 sky130_fd_sc_hd__xnor2_2 _4830_ (.A(_0800_),
    .B(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__a21o_1 _4831_ (.A1(_0730_),
    .A2(_0764_),
    .B1(_0763_),
    .X(_0838_));
 sky130_fd_sc_hd__nand2b_1 _4832_ (.A_N(_0837_),
    .B(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__xnor2_2 _4833_ (.A(_0837_),
    .B(_0838_),
    .Y(_0840_));
 sky130_fd_sc_hd__xnor2_1 _4834_ (.A(_0780_),
    .B(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__a21oi_1 _4835_ (.A1(_0708_),
    .A2(_0768_),
    .B1(_0767_),
    .Y(_0842_));
 sky130_fd_sc_hd__or2_1 _4836_ (.A(_0841_),
    .B(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__xor2_1 _4837_ (.A(_0841_),
    .B(_0842_),
    .X(_0844_));
 sky130_fd_sc_hd__nand2b_1 _4838_ (.A_N(_0706_),
    .B(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__xnor2_1 _4839_ (.A(_0706_),
    .B(_0844_),
    .Y(_0846_));
 sky130_fd_sc_hd__nand2_1 _4840_ (.A(_0772_),
    .B(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__or2_1 _4841_ (.A(_0772_),
    .B(_0846_),
    .X(_0848_));
 sky130_fd_sc_hd__and2_2 _4842_ (.A(_0847_),
    .B(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__a21o_1 _4843_ (.A1(_0691_),
    .A2(_0693_),
    .B1(_0774_),
    .X(_0850_));
 sky130_fd_sc_hd__o31ai_4 _4844_ (.A1(_0696_),
    .A2(_0699_),
    .A3(_0775_),
    .B1(_0850_),
    .Y(_0851_));
 sky130_fd_sc_hd__xnor2_4 _4845_ (.A(_0849_),
    .B(_0851_),
    .Y(_0852_));
 sky130_fd_sc_hd__nand2b_1 _4846_ (.A_N(_0776_),
    .B(_0702_),
    .Y(_0853_));
 sky130_fd_sc_hd__nand2_1 _4847_ (.A(net252),
    .B(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__xor2_2 _4848_ (.A(_0852_),
    .B(_0854_),
    .X(\mul_wb.reg_p[14] ));
 sky130_fd_sc_hd__nand3b_2 _4849_ (.A_N(_0776_),
    .B(_0852_),
    .C(_0702_),
    .Y(_0855_));
 sky130_fd_sc_hd__nand2_1 _4850_ (.A(net252),
    .B(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__a21boi_4 _4851_ (.A1(_0849_),
    .A2(_0851_),
    .B1_N(_0847_),
    .Y(_0857_));
 sky130_fd_sc_hd__a21bo_1 _4852_ (.A1(_0783_),
    .A2(_0786_),
    .B1_N(_0784_),
    .X(_0858_));
 sky130_fd_sc_hd__o21a_2 _4853_ (.A1(_0797_),
    .A2(_0799_),
    .B1(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__or3_1 _4854_ (.A(_0797_),
    .B(_0799_),
    .C(_0858_),
    .X(_0860_));
 sky130_fd_sc_hd__nand2b_1 _4855_ (.A_N(_0859_),
    .B(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__nand2_8 _4856_ (.A(net269),
    .B(net242),
    .Y(_0862_));
 sky130_fd_sc_hd__o21ai_4 _4857_ (.A1(net177),
    .A2(_0862_),
    .B1(_0861_),
    .Y(_0863_));
 sky130_fd_sc_hd__o21ai_4 _4858_ (.A1(_0792_),
    .A2(_0793_),
    .B1(_0795_),
    .Y(_0864_));
 sky130_fd_sc_hd__o21bai_2 _4859_ (.A1(_0802_),
    .A2(_0810_),
    .B1_N(_0809_),
    .Y(_0865_));
 sky130_fd_sc_hd__o22a_1 _4860_ (.A1(net205),
    .A2(net189),
    .B1(net219),
    .B2(_3683_),
    .X(_0866_));
 sky130_fd_sc_hd__or4_1 _4861_ (.A(net208),
    .B(net205),
    .C(net190),
    .D(net219),
    .X(_0867_));
 sky130_fd_sc_hd__and2b_1 _4862_ (.A_N(_0866_),
    .B(_0867_),
    .X(_0868_));
 sky130_fd_sc_hd__nor2_2 _4863_ (.A(net173),
    .B(net217),
    .Y(_0869_));
 sky130_fd_sc_hd__xnor2_4 _4864_ (.A(_0868_),
    .B(_0869_),
    .Y(_0870_));
 sky130_fd_sc_hd__o22a_1 _4865_ (.A1(net197),
    .A2(net192),
    .B1(net223),
    .B2(net201),
    .X(_0871_));
 sky130_fd_sc_hd__or4_1 _4866_ (.A(net201),
    .B(net197),
    .C(net192),
    .D(net223),
    .X(_0872_));
 sky130_fd_sc_hd__and2b_1 _4867_ (.A_N(_0871_),
    .B(_0872_),
    .X(_0873_));
 sky130_fd_sc_hd__nor2_1 _4868_ (.A(net198),
    .B(net191),
    .Y(_0874_));
 sky130_fd_sc_hd__xnor2_1 _4869_ (.A(_0873_),
    .B(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__o31a_1 _4870_ (.A1(net204),
    .A2(net191),
    .A3(_0788_),
    .B1(_0789_),
    .X(_0876_));
 sky130_fd_sc_hd__or2_1 _4871_ (.A(_0875_),
    .B(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__nand2_1 _4872_ (.A(_0875_),
    .B(_0876_),
    .Y(_0878_));
 sky130_fd_sc_hd__nand2_2 _4873_ (.A(_0877_),
    .B(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__xnor2_2 _4874_ (.A(_0870_),
    .B(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__and2b_1 _4875_ (.A_N(_0880_),
    .B(_0865_),
    .X(_0881_));
 sky130_fd_sc_hd__xnor2_2 _4876_ (.A(_0865_),
    .B(_0880_),
    .Y(_0882_));
 sky130_fd_sc_hd__xor2_4 _4877_ (.A(_0864_),
    .B(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__a21bo_1 _4878_ (.A1(_0806_),
    .A2(_0807_),
    .B1_N(_0805_),
    .X(_0884_));
 sky130_fd_sc_hd__o32a_1 _4879_ (.A1(net175),
    .A2(_0815_),
    .A3(net237),
    .B1(_0813_),
    .B2(_0814_),
    .X(_0885_));
 sky130_fd_sc_hd__or2_1 _4880_ (.A(net207),
    .B(_0667_),
    .X(_0886_));
 sky130_fd_sc_hd__a21oi_1 _4881_ (.A1(net212),
    .A2(net211),
    .B1(net237),
    .Y(_0887_));
 sky130_fd_sc_hd__or3_1 _4882_ (.A(_3614_),
    .B(_0816_),
    .C(_0886_),
    .X(_0888_));
 sky130_fd_sc_hd__xnor2_1 _4883_ (.A(_0886_),
    .B(_0887_),
    .Y(_0889_));
 sky130_fd_sc_hd__and3_1 _4884_ (.A(_3526_),
    .B(_3738_),
    .C(_0597_),
    .X(_0890_));
 sky130_fd_sc_hd__xnor2_1 _4885_ (.A(_0889_),
    .B(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__nor2_1 _4886_ (.A(_0885_),
    .B(_0891_),
    .Y(_0892_));
 sky130_fd_sc_hd__xor2_1 _4887_ (.A(_0885_),
    .B(_0891_),
    .X(_0893_));
 sky130_fd_sc_hd__and2_1 _4888_ (.A(_0884_),
    .B(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__nor2_1 _4889_ (.A(_0884_),
    .B(_0893_),
    .Y(_0895_));
 sky130_fd_sc_hd__nor2_2 _4890_ (.A(_0894_),
    .B(_0895_),
    .Y(_0896_));
 sky130_fd_sc_hd__o22ai_1 _4891_ (.A1(net203),
    .A2(net222),
    .B1(_0753_),
    .B2(net209),
    .Y(_0897_));
 sky130_fd_sc_hd__or4_2 _4892_ (.A(net209),
    .B(net203),
    .C(net222),
    .D(_0753_),
    .X(_0898_));
 sky130_fd_sc_hd__nand2_8 _4893_ (.A(net269),
    .B(net247),
    .Y(_0899_));
 sky130_fd_sc_hd__a2bb2o_2 _4894_ (.A1_N(net175),
    .A2_N(_0899_),
    .B1(_0898_),
    .B2(_0897_),
    .X(_0900_));
 sky130_fd_sc_hd__nor2_2 _4895_ (.A(net195),
    .B(net194),
    .Y(_0901_));
 sky130_fd_sc_hd__or2_2 _4896_ (.A(net206),
    .B(net220),
    .X(_0902_));
 sky130_fd_sc_hd__a21oi_2 _4897_ (.A1(_3583_),
    .A2(_3586_),
    .B1(_0822_),
    .Y(_0903_));
 sky130_fd_sc_hd__or3_1 _4898_ (.A(net174),
    .B(_0822_),
    .C(_0902_),
    .X(_0904_));
 sky130_fd_sc_hd__xnor2_4 _4899_ (.A(_0902_),
    .B(_0903_),
    .Y(_0905_));
 sky130_fd_sc_hd__xnor2_4 _4900_ (.A(_0901_),
    .B(_0905_),
    .Y(_0906_));
 sky130_fd_sc_hd__a21oi_2 _4901_ (.A1(_0819_),
    .A2(_0825_),
    .B1(_0824_),
    .Y(_0907_));
 sky130_fd_sc_hd__nor2_1 _4902_ (.A(_0906_),
    .B(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__xor2_4 _4903_ (.A(_0906_),
    .B(_0907_),
    .X(_0909_));
 sky130_fd_sc_hd__xnor2_4 _4904_ (.A(_0900_),
    .B(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__o21ba_2 _4905_ (.A1(_0818_),
    .A2(_0828_),
    .B1_N(_0827_),
    .X(_0911_));
 sky130_fd_sc_hd__nor2_1 _4906_ (.A(_0910_),
    .B(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__xor2_4 _4907_ (.A(_0910_),
    .B(_0911_),
    .X(_0913_));
 sky130_fd_sc_hd__xnor2_4 _4908_ (.A(_0896_),
    .B(_0913_),
    .Y(_0914_));
 sky130_fd_sc_hd__a21bo_2 _4909_ (.A1(_0812_),
    .A2(_0832_),
    .B1_N(_0831_),
    .X(_0915_));
 sky130_fd_sc_hd__nand2b_1 _4910_ (.A_N(_0914_),
    .B(_0915_),
    .Y(_0916_));
 sky130_fd_sc_hd__xnor2_4 _4911_ (.A(_0914_),
    .B(_0915_),
    .Y(_0917_));
 sky130_fd_sc_hd__xnor2_4 _4912_ (.A(_0883_),
    .B(_0917_),
    .Y(_0918_));
 sky130_fd_sc_hd__a21oi_4 _4913_ (.A1(_0800_),
    .A2(_0836_),
    .B1(_0835_),
    .Y(_0919_));
 sky130_fd_sc_hd__nor2_1 _4914_ (.A(_0918_),
    .B(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__xor2_4 _4915_ (.A(_0918_),
    .B(_0919_),
    .X(_0921_));
 sky130_fd_sc_hd__xnor2_2 _4916_ (.A(_0863_),
    .B(_0921_),
    .Y(_0922_));
 sky130_fd_sc_hd__a21boi_2 _4917_ (.A1(_0780_),
    .A2(_0840_),
    .B1_N(_0839_),
    .Y(_0923_));
 sky130_fd_sc_hd__nor2_1 _4918_ (.A(_0922_),
    .B(_0923_),
    .Y(_0924_));
 sky130_fd_sc_hd__xor2_2 _4919_ (.A(_0922_),
    .B(_0923_),
    .X(_0925_));
 sky130_fd_sc_hd__xnor2_1 _4920_ (.A(_0778_),
    .B(_0925_),
    .Y(_0926_));
 sky130_fd_sc_hd__a21oi_1 _4921_ (.A1(_0843_),
    .A2(_0845_),
    .B1(_0926_),
    .Y(_0927_));
 sky130_fd_sc_hd__a21o_1 _4922_ (.A1(_0843_),
    .A2(_0845_),
    .B1(_0926_),
    .X(_0928_));
 sky130_fd_sc_hd__and3_1 _4923_ (.A(_0843_),
    .B(_0845_),
    .C(_0926_),
    .X(_0929_));
 sky130_fd_sc_hd__nor2_2 _4924_ (.A(_0927_),
    .B(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__xnor2_4 _4925_ (.A(_0857_),
    .B(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__xnor2_1 _4926_ (.A(_0856_),
    .B(_0931_),
    .Y(\mul_wb.reg_p[15] ));
 sky130_fd_sc_hd__a21oi_1 _4927_ (.A1(_0864_),
    .A2(_0882_),
    .B1(_0881_),
    .Y(_0932_));
 sky130_fd_sc_hd__o31a_1 _4928_ (.A1(net173),
    .A2(net217),
    .A3(_0866_),
    .B1(_0867_),
    .X(_0933_));
 sky130_fd_sc_hd__nor2_2 _4929_ (.A(_0932_),
    .B(_0933_),
    .Y(_0934_));
 sky130_fd_sc_hd__xnor2_1 _4930_ (.A(_0932_),
    .B(_0933_),
    .Y(_0935_));
 sky130_fd_sc_hd__o21ai_4 _4931_ (.A1(_3587_),
    .A2(_0862_),
    .B1(_0935_),
    .Y(_0936_));
 sky130_fd_sc_hd__o21ai_4 _4932_ (.A1(_0870_),
    .A2(_0879_),
    .B1(_0877_),
    .Y(_0937_));
 sky130_fd_sc_hd__or2_1 _4933_ (.A(_3722_),
    .B(net219),
    .X(_0938_));
 sky130_fd_sc_hd__nor2_1 _4934_ (.A(net198),
    .B(net189),
    .Y(_0939_));
 sky130_fd_sc_hd__xnor2_1 _4935_ (.A(_0938_),
    .B(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__inv_2 _4936_ (.A(_0940_),
    .Y(_0941_));
 sky130_fd_sc_hd__or2_1 _4937_ (.A(net208),
    .B(net217),
    .X(_0942_));
 sky130_fd_sc_hd__xnor2_1 _4938_ (.A(_0940_),
    .B(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__o22ai_1 _4939_ (.A1(net197),
    .A2(net223),
    .B1(net222),
    .B2(net201),
    .Y(_0944_));
 sky130_fd_sc_hd__or4_1 _4940_ (.A(net201),
    .B(net197),
    .C(net223),
    .D(net222),
    .X(_0945_));
 sky130_fd_sc_hd__nand2_1 _4941_ (.A(_0944_),
    .B(_0945_),
    .Y(_0946_));
 sky130_fd_sc_hd__nor2_1 _4942_ (.A(_0346_),
    .B(_0442_),
    .Y(_0947_));
 sky130_fd_sc_hd__xnor2_1 _4943_ (.A(_0946_),
    .B(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__o31a_1 _4944_ (.A1(net199),
    .A2(net191),
    .A3(_0871_),
    .B1(_0872_),
    .X(_0949_));
 sky130_fd_sc_hd__nand2b_1 _4945_ (.A_N(_0949_),
    .B(_0948_),
    .Y(_0950_));
 sky130_fd_sc_hd__xnor2_1 _4946_ (.A(_0948_),
    .B(_0949_),
    .Y(_0951_));
 sky130_fd_sc_hd__xor2_1 _4947_ (.A(_0943_),
    .B(_0951_),
    .X(_0952_));
 sky130_fd_sc_hd__o21a_1 _4948_ (.A1(_0892_),
    .A2(_0894_),
    .B1(_0952_),
    .X(_0953_));
 sky130_fd_sc_hd__nor3_1 _4949_ (.A(_0892_),
    .B(_0894_),
    .C(_0952_),
    .Y(_0954_));
 sky130_fd_sc_hd__nor2_2 _4950_ (.A(_0953_),
    .B(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__xor2_4 _4951_ (.A(_0937_),
    .B(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__a21bo_1 _4952_ (.A1(_0889_),
    .A2(_0890_),
    .B1_N(_0888_),
    .X(_0957_));
 sky130_fd_sc_hd__o22ai_1 _4953_ (.A1(net207),
    .A2(_0753_),
    .B1(_0899_),
    .B2(_3614_),
    .Y(_0958_));
 sky130_fd_sc_hd__and3_1 _4954_ (.A(_3526_),
    .B(_3738_),
    .C(_0668_),
    .X(_0959_));
 sky130_fd_sc_hd__and2_1 _4955_ (.A(_0958_),
    .B(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__xor2_1 _4956_ (.A(_0958_),
    .B(_0959_),
    .X(_0961_));
 sky130_fd_sc_hd__and2b_1 _4957_ (.A_N(_0898_),
    .B(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__xor2_1 _4958_ (.A(_0898_),
    .B(_0961_),
    .X(_0963_));
 sky130_fd_sc_hd__and2b_1 _4959_ (.A_N(_0963_),
    .B(_0957_),
    .X(_0964_));
 sky130_fd_sc_hd__and2b_1 _4960_ (.A_N(_0957_),
    .B(_0963_),
    .X(_0965_));
 sky130_fd_sc_hd__nor2_2 _4961_ (.A(_0964_),
    .B(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__or4_2 _4962_ (.A(net209),
    .B(net203),
    .C(net221),
    .D(_0816_),
    .X(_0967_));
 sky130_fd_sc_hd__o22ai_1 _4963_ (.A1(net203),
    .A2(net221),
    .B1(_0816_),
    .B2(net209),
    .Y(_0968_));
 sky130_fd_sc_hd__and2_2 _4964_ (.A(_0967_),
    .B(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__or2_2 _4965_ (.A(net194),
    .B(net192),
    .X(_0970_));
 sky130_fd_sc_hd__nor2_2 _4966_ (.A(net204),
    .B(net220),
    .Y(_0971_));
 sky130_fd_sc_hd__a21oi_4 _4967_ (.A1(_3648_),
    .A2(_3656_),
    .B1(_0822_),
    .Y(_0972_));
 sky130_fd_sc_hd__nand2_1 _4968_ (.A(_0971_),
    .B(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__xnor2_4 _4969_ (.A(_0971_),
    .B(_0972_),
    .Y(_0974_));
 sky130_fd_sc_hd__xnor2_4 _4970_ (.A(_0970_),
    .B(_0974_),
    .Y(_0975_));
 sky130_fd_sc_hd__a21boi_4 _4971_ (.A1(_0901_),
    .A2(_0905_),
    .B1_N(_0904_),
    .Y(_0976_));
 sky130_fd_sc_hd__nor2_1 _4972_ (.A(_0975_),
    .B(_0976_),
    .Y(_0977_));
 sky130_fd_sc_hd__xor2_4 _4973_ (.A(_0975_),
    .B(_0976_),
    .X(_0978_));
 sky130_fd_sc_hd__xnor2_4 _4974_ (.A(_0969_),
    .B(_0978_),
    .Y(_0979_));
 sky130_fd_sc_hd__a21oi_4 _4975_ (.A1(_0900_),
    .A2(_0909_),
    .B1(_0908_),
    .Y(_0980_));
 sky130_fd_sc_hd__nor2_1 _4976_ (.A(_0979_),
    .B(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__xor2_4 _4977_ (.A(_0979_),
    .B(_0980_),
    .X(_0982_));
 sky130_fd_sc_hd__xnor2_4 _4978_ (.A(_0966_),
    .B(_0982_),
    .Y(_0983_));
 sky130_fd_sc_hd__a21o_2 _4979_ (.A1(_0896_),
    .A2(_0913_),
    .B1(_0912_),
    .X(_0984_));
 sky130_fd_sc_hd__and2b_1 _4980_ (.A_N(_0983_),
    .B(_0984_),
    .X(_0985_));
 sky130_fd_sc_hd__xnor2_4 _4981_ (.A(_0983_),
    .B(_0984_),
    .Y(_0986_));
 sky130_fd_sc_hd__xnor2_4 _4982_ (.A(_0956_),
    .B(_0986_),
    .Y(_0987_));
 sky130_fd_sc_hd__a21boi_4 _4983_ (.A1(_0883_),
    .A2(_0917_),
    .B1_N(_0916_),
    .Y(_0988_));
 sky130_fd_sc_hd__nor2_1 _4984_ (.A(_0987_),
    .B(_0988_),
    .Y(_0989_));
 sky130_fd_sc_hd__xor2_4 _4985_ (.A(_0987_),
    .B(_0988_),
    .X(_0990_));
 sky130_fd_sc_hd__xnor2_4 _4986_ (.A(_0936_),
    .B(_0990_),
    .Y(_0991_));
 sky130_fd_sc_hd__a21oi_4 _4987_ (.A1(_0863_),
    .A2(_0921_),
    .B1(_0920_),
    .Y(_0992_));
 sky130_fd_sc_hd__nor2_1 _4988_ (.A(_0991_),
    .B(_0992_),
    .Y(_0993_));
 sky130_fd_sc_hd__xor2_4 _4989_ (.A(_0991_),
    .B(_0992_),
    .X(_0994_));
 sky130_fd_sc_hd__xnor2_4 _4990_ (.A(_0859_),
    .B(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__a21oi_4 _4991_ (.A1(_0778_),
    .A2(_0925_),
    .B1(_0924_),
    .Y(_0996_));
 sky130_fd_sc_hd__nor2_1 _4992_ (.A(_0995_),
    .B(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__xor2_4 _4993_ (.A(_0995_),
    .B(_0996_),
    .X(_0998_));
 sky130_fd_sc_hd__a21oi_1 _4994_ (.A1(_0847_),
    .A2(_0928_),
    .B1(_0929_),
    .Y(_0999_));
 sky130_fd_sc_hd__a31o_4 _4995_ (.A1(_0849_),
    .A2(_0851_),
    .A3(_0930_),
    .B1(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__xnor2_4 _4996_ (.A(_0998_),
    .B(_1000_),
    .Y(_1001_));
 sky130_fd_sc_hd__nor2_1 _4997_ (.A(_0855_),
    .B(_0931_),
    .Y(_1002_));
 sky130_fd_sc_hd__nor2_1 _4998_ (.A(_3620_),
    .B(_1002_),
    .Y(_1003_));
 sky130_fd_sc_hd__xnor2_1 _4999_ (.A(_1001_),
    .B(_1003_),
    .Y(\mul_wb.reg_p[16] ));
 sky130_fd_sc_hd__a21oi_1 _5000_ (.A1(_1001_),
    .A2(_1002_),
    .B1(_3620_),
    .Y(_1004_));
 sky130_fd_sc_hd__a21o_1 _5001_ (.A1(_0998_),
    .A2(_1000_),
    .B1(_0997_),
    .X(_1005_));
 sky130_fd_sc_hd__a21oi_1 _5002_ (.A1(_0937_),
    .A2(_0955_),
    .B1(_0953_),
    .Y(_1006_));
 sky130_fd_sc_hd__o32a_1 _5003_ (.A1(net199),
    .A2(net189),
    .A3(_0938_),
    .B1(_0941_),
    .B2(_0942_),
    .X(_1007_));
 sky130_fd_sc_hd__or2_4 _5004_ (.A(_1006_),
    .B(_1007_),
    .X(_1008_));
 sky130_fd_sc_hd__nand2_1 _5005_ (.A(_1006_),
    .B(_1007_),
    .Y(_1009_));
 sky130_fd_sc_hd__a2bb2o_2 _5006_ (.A1_N(net173),
    .A2_N(_0862_),
    .B1(_1008_),
    .B2(_1009_),
    .X(_1010_));
 sky130_fd_sc_hd__a21bo_2 _5007_ (.A1(_0943_),
    .A2(_0951_),
    .B1_N(_0950_),
    .X(_1011_));
 sky130_fd_sc_hd__o22a_1 _5008_ (.A1(_0346_),
    .A2(net190),
    .B1(net219),
    .B2(net205),
    .X(_1012_));
 sky130_fd_sc_hd__or4_1 _5009_ (.A(net205),
    .B(_0346_),
    .C(net190),
    .D(net219),
    .X(_1013_));
 sky130_fd_sc_hd__and2b_1 _5010_ (.A_N(_1012_),
    .B(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__or2_1 _5011_ (.A(_3722_),
    .B(net217),
    .X(_1015_));
 sky130_fd_sc_hd__xor2_2 _5012_ (.A(_1014_),
    .B(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__o22a_1 _5013_ (.A1(net197),
    .A2(_0535_),
    .B1(_0598_),
    .B2(net200),
    .X(_1017_));
 sky130_fd_sc_hd__or4_1 _5014_ (.A(net201),
    .B(net197),
    .C(_0535_),
    .D(_0598_),
    .X(_1018_));
 sky130_fd_sc_hd__nand2b_1 _5015_ (.A_N(_1017_),
    .B(_1018_),
    .Y(_1019_));
 sky130_fd_sc_hd__nor2_1 _5016_ (.A(net193),
    .B(_0442_),
    .Y(_1020_));
 sky130_fd_sc_hd__xnor2_2 _5017_ (.A(_1019_),
    .B(_1020_),
    .Y(_1021_));
 sky130_fd_sc_hd__a21bo_1 _5018_ (.A1(_0944_),
    .A2(_0947_),
    .B1_N(_0945_),
    .X(_1022_));
 sky130_fd_sc_hd__nand2_1 _5019_ (.A(_1021_),
    .B(_1022_),
    .Y(_1023_));
 sky130_fd_sc_hd__nor2_1 _5020_ (.A(_1021_),
    .B(_1022_),
    .Y(_1024_));
 sky130_fd_sc_hd__xor2_1 _5021_ (.A(_1021_),
    .B(_1022_),
    .X(_1025_));
 sky130_fd_sc_hd__xnor2_1 _5022_ (.A(_1016_),
    .B(_1025_),
    .Y(_1026_));
 sky130_fd_sc_hd__o21a_1 _5023_ (.A1(_0962_),
    .A2(_0964_),
    .B1(_1026_),
    .X(_1027_));
 sky130_fd_sc_hd__nor3_1 _5024_ (.A(_0962_),
    .B(_0964_),
    .C(_1026_),
    .Y(_1028_));
 sky130_fd_sc_hd__or2_2 _5025_ (.A(_1027_),
    .B(_1028_),
    .X(_1029_));
 sky130_fd_sc_hd__and2b_1 _5026_ (.A_N(_1029_),
    .B(_1011_),
    .X(_1030_));
 sky130_fd_sc_hd__xnor2_4 _5027_ (.A(_1011_),
    .B(_1029_),
    .Y(_1031_));
 sky130_fd_sc_hd__nor2_1 _5028_ (.A(net207),
    .B(_0816_),
    .Y(_1032_));
 sky130_fd_sc_hd__or2_1 _5029_ (.A(net207),
    .B(net237),
    .X(_1033_));
 sky130_fd_sc_hd__and4_2 _5030_ (.A(_3526_),
    .B(_3738_),
    .C(_0752_),
    .D(_1032_),
    .X(_1034_));
 sky130_fd_sc_hd__a31oi_2 _5031_ (.A1(_3526_),
    .A2(_3738_),
    .A3(_0752_),
    .B1(_1032_),
    .Y(_1035_));
 sky130_fd_sc_hd__nor3_1 _5032_ (.A(_0967_),
    .B(_1034_),
    .C(_1035_),
    .Y(_1036_));
 sky130_fd_sc_hd__or3_1 _5033_ (.A(_0967_),
    .B(_1034_),
    .C(_1035_),
    .X(_1037_));
 sky130_fd_sc_hd__o21ai_1 _5034_ (.A1(_1034_),
    .A2(_1035_),
    .B1(_0967_),
    .Y(_1038_));
 sky130_fd_sc_hd__and3_1 _5035_ (.A(_0960_),
    .B(_1037_),
    .C(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__a21oi_1 _5036_ (.A1(_1037_),
    .A2(_1038_),
    .B1(_0960_),
    .Y(_1040_));
 sky130_fd_sc_hd__or2_2 _5037_ (.A(_1039_),
    .B(_1040_),
    .X(_1041_));
 sky130_fd_sc_hd__inv_2 _5038_ (.A(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__o22a_2 _5039_ (.A1(net203),
    .A2(net227),
    .B1(_0899_),
    .B2(net209),
    .X(_1043_));
 sky130_fd_sc_hd__nor2_2 _5040_ (.A(net194),
    .B(net223),
    .Y(_1044_));
 sky130_fd_sc_hd__o22a_1 _5041_ (.A1(net199),
    .A2(net220),
    .B1(_0822_),
    .B2(net208),
    .X(_1045_));
 sky130_fd_sc_hd__or4_1 _5042_ (.A(net208),
    .B(net198),
    .C(net220),
    .D(_0822_),
    .X(_1046_));
 sky130_fd_sc_hd__and2b_1 _5043_ (.A_N(_1045_),
    .B(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__xnor2_4 _5044_ (.A(_1044_),
    .B(_1047_),
    .Y(_1048_));
 sky130_fd_sc_hd__o31a_2 _5045_ (.A1(net194),
    .A2(net192),
    .A3(_0974_),
    .B1(_0973_),
    .X(_1049_));
 sky130_fd_sc_hd__or2_1 _5046_ (.A(_1048_),
    .B(_1049_),
    .X(_1050_));
 sky130_fd_sc_hd__xnor2_4 _5047_ (.A(_1048_),
    .B(_1049_),
    .Y(_1051_));
 sky130_fd_sc_hd__xnor2_4 _5048_ (.A(_1043_),
    .B(_1051_),
    .Y(_1052_));
 sky130_fd_sc_hd__a21oi_4 _5049_ (.A1(_0969_),
    .A2(_0978_),
    .B1(_0977_),
    .Y(_1053_));
 sky130_fd_sc_hd__nor2_1 _5050_ (.A(_1052_),
    .B(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__xor2_4 _5051_ (.A(_1052_),
    .B(_1053_),
    .X(_1055_));
 sky130_fd_sc_hd__xnor2_4 _5052_ (.A(_1041_),
    .B(_1055_),
    .Y(_1056_));
 sky130_fd_sc_hd__a21oi_2 _5053_ (.A1(_0966_),
    .A2(_0982_),
    .B1(_0981_),
    .Y(_1057_));
 sky130_fd_sc_hd__and2b_1 _5054_ (.A_N(_1057_),
    .B(_1056_),
    .X(_1058_));
 sky130_fd_sc_hd__xnor2_4 _5055_ (.A(_1056_),
    .B(_1057_),
    .Y(_1059_));
 sky130_fd_sc_hd__xnor2_4 _5056_ (.A(_1031_),
    .B(_1059_),
    .Y(_1060_));
 sky130_fd_sc_hd__a21oi_4 _5057_ (.A1(_0956_),
    .A2(_0986_),
    .B1(_0985_),
    .Y(_1061_));
 sky130_fd_sc_hd__nor2_1 _5058_ (.A(_1060_),
    .B(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__xor2_4 _5059_ (.A(_1060_),
    .B(_1061_),
    .X(_1063_));
 sky130_fd_sc_hd__xnor2_4 _5060_ (.A(_1010_),
    .B(_1063_),
    .Y(_1064_));
 sky130_fd_sc_hd__a21oi_2 _5061_ (.A1(_0936_),
    .A2(_0990_),
    .B1(_0989_),
    .Y(_1065_));
 sky130_fd_sc_hd__nor2_1 _5062_ (.A(_1064_),
    .B(_1065_),
    .Y(_1066_));
 sky130_fd_sc_hd__xor2_4 _5063_ (.A(_1064_),
    .B(_1065_),
    .X(_1067_));
 sky130_fd_sc_hd__xnor2_4 _5064_ (.A(_0934_),
    .B(_1067_),
    .Y(_1068_));
 sky130_fd_sc_hd__a21oi_4 _5065_ (.A1(_0859_),
    .A2(_0994_),
    .B1(_0993_),
    .Y(_1069_));
 sky130_fd_sc_hd__and2_1 _5066_ (.A(_1068_),
    .B(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__xor2_4 _5067_ (.A(_1068_),
    .B(_1069_),
    .X(_1071_));
 sky130_fd_sc_hd__xnor2_4 _5068_ (.A(_1005_),
    .B(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__xnor2_1 _5069_ (.A(_1004_),
    .B(_1072_),
    .Y(\mul_wb.reg_p[17] ));
 sky130_fd_sc_hd__o21ai_1 _5070_ (.A1(_1012_),
    .A2(_1015_),
    .B1(_1013_),
    .Y(_1073_));
 sky130_fd_sc_hd__o21a_2 _5071_ (.A1(_1027_),
    .A2(_1030_),
    .B1(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__nor3_1 _5072_ (.A(_1027_),
    .B(_1030_),
    .C(_1073_),
    .Y(_1075_));
 sky130_fd_sc_hd__o22ai_4 _5073_ (.A1(net208),
    .A2(_0862_),
    .B1(_1074_),
    .B2(_1075_),
    .Y(_1076_));
 sky130_fd_sc_hd__o21ai_4 _5074_ (.A1(_1016_),
    .A2(_1024_),
    .B1(_1023_),
    .Y(_1077_));
 sky130_fd_sc_hd__o22ai_1 _5075_ (.A1(net193),
    .A2(net189),
    .B1(net219),
    .B2(net199),
    .Y(_1078_));
 sky130_fd_sc_hd__or4_1 _5076_ (.A(net199),
    .B(net193),
    .C(net189),
    .D(net219),
    .X(_1079_));
 sky130_fd_sc_hd__nand2_1 _5077_ (.A(_1078_),
    .B(_1079_),
    .Y(_1080_));
 sky130_fd_sc_hd__nor2_1 _5078_ (.A(net205),
    .B(_0715_),
    .Y(_1081_));
 sky130_fd_sc_hd__xnor2_1 _5079_ (.A(_1080_),
    .B(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__o22ai_2 _5080_ (.A1(net197),
    .A2(net221),
    .B1(net227),
    .B2(net201),
    .Y(_1083_));
 sky130_fd_sc_hd__or4_1 _5081_ (.A(net201),
    .B(net197),
    .C(_0598_),
    .D(net227),
    .X(_1084_));
 sky130_fd_sc_hd__nand2_1 _5082_ (.A(_1083_),
    .B(_1084_),
    .Y(_1085_));
 sky130_fd_sc_hd__nor2_1 _5083_ (.A(_0442_),
    .B(net224),
    .Y(_1086_));
 sky130_fd_sc_hd__xnor2_1 _5084_ (.A(_1085_),
    .B(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__o31ai_2 _5085_ (.A1(net193),
    .A2(_0442_),
    .A3(_1017_),
    .B1(_1018_),
    .Y(_1088_));
 sky130_fd_sc_hd__nand2_1 _5086_ (.A(_1087_),
    .B(_1088_),
    .Y(_1089_));
 sky130_fd_sc_hd__xor2_1 _5087_ (.A(_1087_),
    .B(_1088_),
    .X(_1090_));
 sky130_fd_sc_hd__nand2_1 _5088_ (.A(_1082_),
    .B(_1090_),
    .Y(_1091_));
 sky130_fd_sc_hd__xnor2_1 _5089_ (.A(_1082_),
    .B(_1090_),
    .Y(_1092_));
 sky130_fd_sc_hd__o21ba_1 _5090_ (.A1(_1036_),
    .A2(_1039_),
    .B1_N(_1092_),
    .X(_1093_));
 sky130_fd_sc_hd__or3b_1 _5091_ (.A(_1036_),
    .B(_1039_),
    .C_N(_1092_),
    .X(_1094_));
 sky130_fd_sc_hd__and2b_2 _5092_ (.A_N(_1093_),
    .B(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__xor2_4 _5093_ (.A(_1077_),
    .B(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__o22a_1 _5094_ (.A1(_3739_),
    .A2(_0816_),
    .B1(_0899_),
    .B2(_3697_),
    .X(_1097_));
 sky130_fd_sc_hd__nor2_2 _5095_ (.A(_1034_),
    .B(_1097_),
    .Y(_1098_));
 sky130_fd_sc_hd__nor2_1 _5096_ (.A(net194),
    .B(net222),
    .Y(_1099_));
 sky130_fd_sc_hd__a31o_1 _5097_ (.A1(_3717_),
    .A2(_3718_),
    .A3(_3721_),
    .B1(_0822_),
    .X(_1100_));
 sky130_fd_sc_hd__o211a_1 _5098_ (.A1(_0341_),
    .A2(_0345_),
    .B1(_0606_),
    .C1(_3415_),
    .X(_1101_));
 sky130_fd_sc_hd__or3_1 _5099_ (.A(net195),
    .B(net220),
    .C(_1100_),
    .X(_1102_));
 sky130_fd_sc_hd__xnor2_1 _5100_ (.A(_1100_),
    .B(_1101_),
    .Y(_1103_));
 sky130_fd_sc_hd__xnor2_1 _5101_ (.A(_1099_),
    .B(_1103_),
    .Y(_1104_));
 sky130_fd_sc_hd__o31a_1 _5102_ (.A1(net194),
    .A2(net223),
    .A3(_1045_),
    .B1(_1046_),
    .X(_1105_));
 sky130_fd_sc_hd__nor2_1 _5103_ (.A(_1104_),
    .B(_1105_),
    .Y(_1106_));
 sky130_fd_sc_hd__xnor2_1 _5104_ (.A(_1104_),
    .B(_1105_),
    .Y(_1107_));
 sky130_fd_sc_hd__nor3_2 _5105_ (.A(net203),
    .B(_0753_),
    .C(_1107_),
    .Y(_1108_));
 sky130_fd_sc_hd__o21a_1 _5106_ (.A1(net203),
    .A2(_0753_),
    .B1(_1107_),
    .X(_1109_));
 sky130_fd_sc_hd__nor2_2 _5107_ (.A(_1108_),
    .B(_1109_),
    .Y(_1110_));
 sky130_fd_sc_hd__o21a_2 _5108_ (.A1(_1043_),
    .A2(_1051_),
    .B1(_1050_),
    .X(_1111_));
 sky130_fd_sc_hd__and2b_1 _5109_ (.A_N(_1111_),
    .B(_1110_),
    .X(_1112_));
 sky130_fd_sc_hd__xnor2_4 _5110_ (.A(_1110_),
    .B(_1111_),
    .Y(_1113_));
 sky130_fd_sc_hd__xor2_4 _5111_ (.A(_1098_),
    .B(_1113_),
    .X(_1114_));
 sky130_fd_sc_hd__a21oi_2 _5112_ (.A1(_1042_),
    .A2(_1055_),
    .B1(_1054_),
    .Y(_1115_));
 sky130_fd_sc_hd__and2b_1 _5113_ (.A_N(_1115_),
    .B(_1114_),
    .X(_1116_));
 sky130_fd_sc_hd__xnor2_4 _5114_ (.A(_1114_),
    .B(_1115_),
    .Y(_1117_));
 sky130_fd_sc_hd__xnor2_4 _5115_ (.A(_1096_),
    .B(_1117_),
    .Y(_1118_));
 sky130_fd_sc_hd__a21oi_2 _5116_ (.A1(_1031_),
    .A2(_1059_),
    .B1(_1058_),
    .Y(_1119_));
 sky130_fd_sc_hd__nor2_1 _5117_ (.A(_1118_),
    .B(_1119_),
    .Y(_1120_));
 sky130_fd_sc_hd__xor2_4 _5118_ (.A(_1118_),
    .B(_1119_),
    .X(_1121_));
 sky130_fd_sc_hd__xnor2_4 _5119_ (.A(_1076_),
    .B(_1121_),
    .Y(_1122_));
 sky130_fd_sc_hd__a21oi_2 _5120_ (.A1(_1010_),
    .A2(_1063_),
    .B1(_1062_),
    .Y(_1123_));
 sky130_fd_sc_hd__or2_1 _5121_ (.A(_1122_),
    .B(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__xnor2_4 _5122_ (.A(_1122_),
    .B(_1123_),
    .Y(_1125_));
 sky130_fd_sc_hd__xnor2_4 _5123_ (.A(_1008_),
    .B(_1125_),
    .Y(_1126_));
 sky130_fd_sc_hd__a21oi_4 _5124_ (.A1(_0934_),
    .A2(_1067_),
    .B1(_1066_),
    .Y(_1127_));
 sky130_fd_sc_hd__or2_1 _5125_ (.A(_1126_),
    .B(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__xnor2_4 _5126_ (.A(_1126_),
    .B(_1127_),
    .Y(_1129_));
 sky130_fd_sc_hd__o22a_1 _5127_ (.A1(_0995_),
    .A2(_0996_),
    .B1(_1068_),
    .B2(_1069_),
    .X(_1130_));
 sky130_fd_sc_hd__and2_1 _5128_ (.A(_0998_),
    .B(_1071_),
    .X(_1131_));
 sky130_fd_sc_hd__o2bb2a_2 _5129_ (.A1_N(_1000_),
    .A2_N(_1131_),
    .B1(_1130_),
    .B2(_1070_),
    .X(_1132_));
 sky130_fd_sc_hd__xnor2_4 _5130_ (.A(_1129_),
    .B(_1132_),
    .Y(_1133_));
 sky130_fd_sc_hd__a31o_1 _5131_ (.A1(_1001_),
    .A2(_1002_),
    .A3(_1072_),
    .B1(_3620_),
    .X(_1134_));
 sky130_fd_sc_hd__xor2_1 _5132_ (.A(_1133_),
    .B(_1134_),
    .X(\mul_wb.reg_p[18] ));
 sky130_fd_sc_hd__nand4_2 _5133_ (.A(_1001_),
    .B(_1002_),
    .C(_1072_),
    .D(_1133_),
    .Y(_1135_));
 sky130_fd_sc_hd__nand2_1 _5134_ (.A(net252),
    .B(_1135_),
    .Y(_1136_));
 sky130_fd_sc_hd__o21ai_4 _5135_ (.A1(_1008_),
    .A2(_1125_),
    .B1(_1124_),
    .Y(_1137_));
 sky130_fd_sc_hd__a21o_1 _5136_ (.A1(_1077_),
    .A2(_1095_),
    .B1(_1093_),
    .X(_1138_));
 sky130_fd_sc_hd__a21bo_1 _5137_ (.A1(_1078_),
    .A2(_1081_),
    .B1_N(_1079_),
    .X(_1139_));
 sky130_fd_sc_hd__nand2_1 _5138_ (.A(_1138_),
    .B(_1139_),
    .Y(_1140_));
 sky130_fd_sc_hd__or2_1 _5139_ (.A(_1138_),
    .B(_1139_),
    .X(_1141_));
 sky130_fd_sc_hd__a2bb2o_1 _5140_ (.A1_N(_3722_),
    .A2_N(_0862_),
    .B1(_1140_),
    .B2(_1141_),
    .X(_1142_));
 sky130_fd_sc_hd__o22ai_1 _5141_ (.A1(net224),
    .A2(net190),
    .B1(net218),
    .B2(net195),
    .Y(_1143_));
 sky130_fd_sc_hd__or4_2 _5142_ (.A(_0346_),
    .B(net224),
    .C(net190),
    .D(net218),
    .X(_1144_));
 sky130_fd_sc_hd__nand2_1 _5143_ (.A(_1143_),
    .B(_1144_),
    .Y(_1145_));
 sky130_fd_sc_hd__nor2_1 _5144_ (.A(net199),
    .B(_0715_),
    .Y(_1146_));
 sky130_fd_sc_hd__or3_2 _5145_ (.A(net199),
    .B(_0715_),
    .C(_1145_),
    .X(_1147_));
 sky130_fd_sc_hd__xnor2_1 _5146_ (.A(_1145_),
    .B(_1146_),
    .Y(_1148_));
 sky130_fd_sc_hd__o211a_1 _5147_ (.A1(_0328_),
    .A2(_0331_),
    .B1(_0668_),
    .C1(_3511_),
    .X(_1149_));
 sky130_fd_sc_hd__o311a_1 _5148_ (.A1(_0265_),
    .A2(_0266_),
    .A3(_0271_),
    .B1(_0752_),
    .C1(_3515_),
    .X(_1150_));
 sky130_fd_sc_hd__xnor2_2 _5149_ (.A(_1149_),
    .B(_1150_),
    .Y(_1151_));
 sky130_fd_sc_hd__nor2_1 _5150_ (.A(net191),
    .B(_0535_),
    .Y(_1152_));
 sky130_fd_sc_hd__o21a_1 _5151_ (.A1(net191),
    .A2(net222),
    .B1(_1151_),
    .X(_1153_));
 sky130_fd_sc_hd__or3_1 _5152_ (.A(net191),
    .B(net222),
    .C(_1151_),
    .X(_1154_));
 sky130_fd_sc_hd__inv_2 _5153_ (.A(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__xnor2_1 _5154_ (.A(_1151_),
    .B(_1152_),
    .Y(_1156_));
 sky130_fd_sc_hd__a21boi_2 _5155_ (.A1(_1083_),
    .A2(_1086_),
    .B1_N(_1084_),
    .Y(_1157_));
 sky130_fd_sc_hd__xnor2_1 _5156_ (.A(_1156_),
    .B(_1157_),
    .Y(_1158_));
 sky130_fd_sc_hd__nand2_1 _5157_ (.A(_1148_),
    .B(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__or2_1 _5158_ (.A(_1148_),
    .B(_1158_),
    .X(_1160_));
 sky130_fd_sc_hd__nand2_1 _5159_ (.A(_1159_),
    .B(_1160_),
    .Y(_1161_));
 sky130_fd_sc_hd__xor2_1 _5160_ (.A(_1034_),
    .B(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__a21o_1 _5161_ (.A1(_1089_),
    .A2(_1091_),
    .B1(_1162_),
    .X(_1163_));
 sky130_fd_sc_hd__nand3_1 _5162_ (.A(_1089_),
    .B(_1091_),
    .C(_1162_),
    .Y(_1164_));
 sky130_fd_sc_hd__nand2_1 _5163_ (.A(_1163_),
    .B(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__nor2_1 _5164_ (.A(net203),
    .B(_0816_),
    .Y(_1166_));
 sky130_fd_sc_hd__or2_1 _5165_ (.A(net194),
    .B(net221),
    .X(_1167_));
 sky130_fd_sc_hd__o311a_1 _5166_ (.A1(_3765_),
    .A2(_3766_),
    .A3(_3772_),
    .B1(_0821_),
    .C1(_3429_),
    .X(_1168_));
 sky130_fd_sc_hd__a311o_1 _5167_ (.A1(_0393_),
    .A2(_0395_),
    .A3(_0398_),
    .B1(net220),
    .C1(_3409_),
    .X(_1169_));
 sky130_fd_sc_hd__or3_1 _5168_ (.A(net205),
    .B(_0822_),
    .C(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__xor2_1 _5169_ (.A(_1168_),
    .B(_1169_),
    .X(_1171_));
 sky130_fd_sc_hd__or2_1 _5170_ (.A(_1167_),
    .B(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__xnor2_1 _5171_ (.A(_1167_),
    .B(_1171_),
    .Y(_1173_));
 sky130_fd_sc_hd__a21bo_1 _5172_ (.A1(_1099_),
    .A2(_1103_),
    .B1_N(_1102_),
    .X(_1174_));
 sky130_fd_sc_hd__and2b_1 _5173_ (.A_N(_1173_),
    .B(_1174_),
    .X(_1175_));
 sky130_fd_sc_hd__nand2b_1 _5174_ (.A_N(_1174_),
    .B(_1173_),
    .Y(_1176_));
 sky130_fd_sc_hd__xor2_1 _5175_ (.A(_1173_),
    .B(_1174_),
    .X(_1177_));
 sky130_fd_sc_hd__xnor2_1 _5176_ (.A(_1166_),
    .B(_1177_),
    .Y(_1178_));
 sky130_fd_sc_hd__o21a_1 _5177_ (.A1(_1106_),
    .A2(_1108_),
    .B1(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__nor3_1 _5178_ (.A(_1106_),
    .B(_1108_),
    .C(_1178_),
    .Y(_1180_));
 sky130_fd_sc_hd__o22a_1 _5179_ (.A1(_3739_),
    .A2(_0899_),
    .B1(_1179_),
    .B2(_1180_),
    .X(_1181_));
 sky130_fd_sc_hd__a21oi_2 _5180_ (.A1(_1098_),
    .A2(_1113_),
    .B1(_1112_),
    .Y(_1182_));
 sky130_fd_sc_hd__or2_1 _5181_ (.A(_1181_),
    .B(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__xnor2_2 _5182_ (.A(_1181_),
    .B(_1182_),
    .Y(_1184_));
 sky130_fd_sc_hd__xnor2_2 _5183_ (.A(_1165_),
    .B(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__a21oi_2 _5184_ (.A1(_1096_),
    .A2(_1117_),
    .B1(_1116_),
    .Y(_1186_));
 sky130_fd_sc_hd__nor2_1 _5185_ (.A(_1185_),
    .B(_1186_),
    .Y(_1187_));
 sky130_fd_sc_hd__xor2_2 _5186_ (.A(_1185_),
    .B(_1186_),
    .X(_1188_));
 sky130_fd_sc_hd__xnor2_2 _5187_ (.A(_1142_),
    .B(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__a21oi_2 _5188_ (.A1(_1076_),
    .A2(_1121_),
    .B1(_1120_),
    .Y(_1190_));
 sky130_fd_sc_hd__nor2_1 _5189_ (.A(_1189_),
    .B(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__nand2_1 _5190_ (.A(_1189_),
    .B(_1190_),
    .Y(_1192_));
 sky130_fd_sc_hd__xnor2_2 _5191_ (.A(_1189_),
    .B(_1190_),
    .Y(_1193_));
 sky130_fd_sc_hd__xnor2_4 _5192_ (.A(_1074_),
    .B(_1193_),
    .Y(_1194_));
 sky130_fd_sc_hd__nand2_1 _5193_ (.A(_1137_),
    .B(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__nor2_1 _5194_ (.A(_1137_),
    .B(_1194_),
    .Y(_1196_));
 sky130_fd_sc_hd__xnor2_4 _5195_ (.A(_1137_),
    .B(_1194_),
    .Y(_1197_));
 sky130_fd_sc_hd__o21ai_2 _5196_ (.A1(_1129_),
    .A2(_1132_),
    .B1(_1128_),
    .Y(_1198_));
 sky130_fd_sc_hd__xnor2_4 _5197_ (.A(_1197_),
    .B(_1198_),
    .Y(_1199_));
 sky130_fd_sc_hd__xnor2_1 _5198_ (.A(_1136_),
    .B(_1199_),
    .Y(\mul_wb.reg_p[19] ));
 sky130_fd_sc_hd__o41a_1 _5199_ (.A1(_3739_),
    .A2(net216),
    .A3(_1033_),
    .A4(_1161_),
    .B1(_1163_),
    .X(_1200_));
 sky130_fd_sc_hd__a21oi_4 _5200_ (.A1(_1144_),
    .A2(_1147_),
    .B1(_1200_),
    .Y(_1201_));
 sky130_fd_sc_hd__and3_1 _5201_ (.A(_1144_),
    .B(_1147_),
    .C(_1200_),
    .X(_1202_));
 sky130_fd_sc_hd__o22ai_4 _5202_ (.A1(net205),
    .A2(_0862_),
    .B1(_1201_),
    .B2(_1202_),
    .Y(_1203_));
 sky130_fd_sc_hd__o31ai_2 _5203_ (.A1(_1153_),
    .A2(_1155_),
    .A3(_1157_),
    .B1(_1159_),
    .Y(_1204_));
 sky130_fd_sc_hd__o22ai_1 _5204_ (.A1(net189),
    .A2(_0535_),
    .B1(net218),
    .B2(net193),
    .Y(_1205_));
 sky130_fd_sc_hd__or4_1 _5205_ (.A(net193),
    .B(net189),
    .C(_0535_),
    .D(net218),
    .X(_1206_));
 sky130_fd_sc_hd__nand2_1 _5206_ (.A(_1205_),
    .B(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__nor2_1 _5207_ (.A(_0346_),
    .B(net217),
    .Y(_1208_));
 sky130_fd_sc_hd__xnor2_1 _5208_ (.A(_1207_),
    .B(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__o22ai_2 _5209_ (.A1(net197),
    .A2(net216),
    .B1(net237),
    .B2(net201),
    .Y(_1210_));
 sky130_fd_sc_hd__or4_1 _5210_ (.A(net201),
    .B(net197),
    .C(net216),
    .D(net237),
    .X(_1211_));
 sky130_fd_sc_hd__nand2_1 _5211_ (.A(_1210_),
    .B(_1211_),
    .Y(_1212_));
 sky130_fd_sc_hd__nor2_1 _5212_ (.A(net191),
    .B(net221),
    .Y(_1213_));
 sky130_fd_sc_hd__xnor2_1 _5213_ (.A(_1212_),
    .B(_1213_),
    .Y(_1214_));
 sky130_fd_sc_hd__a21bo_1 _5214_ (.A1(_1149_),
    .A2(_1150_),
    .B1_N(_1154_),
    .X(_1215_));
 sky130_fd_sc_hd__nand2_1 _5215_ (.A(_1214_),
    .B(_1215_),
    .Y(_1216_));
 sky130_fd_sc_hd__xor2_1 _5216_ (.A(_1214_),
    .B(_1215_),
    .X(_1217_));
 sky130_fd_sc_hd__xnor2_1 _5217_ (.A(_1209_),
    .B(_1217_),
    .Y(_1218_));
 sky130_fd_sc_hd__nand2b_1 _5218_ (.A_N(_1218_),
    .B(_1204_),
    .Y(_1219_));
 sky130_fd_sc_hd__xnor2_1 _5219_ (.A(_1204_),
    .B(_1218_),
    .Y(_1220_));
 sky130_fd_sc_hd__or2_1 _5220_ (.A(net194),
    .B(net227),
    .X(_1221_));
 sky130_fd_sc_hd__o211a_1 _5221_ (.A1(_0281_),
    .A2(_0285_),
    .B1(_0821_),
    .C1(_3417_),
    .X(_1222_));
 sky130_fd_sc_hd__nor2_1 _5222_ (.A(net223),
    .B(net220),
    .Y(_1223_));
 sky130_fd_sc_hd__nand2_1 _5223_ (.A(_1222_),
    .B(_1223_),
    .Y(_1224_));
 sky130_fd_sc_hd__xnor2_1 _5224_ (.A(_1222_),
    .B(_1223_),
    .Y(_1225_));
 sky130_fd_sc_hd__xnor2_1 _5225_ (.A(_1221_),
    .B(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__a21o_1 _5226_ (.A1(_1170_),
    .A2(_1172_),
    .B1(_1226_),
    .X(_1227_));
 sky130_fd_sc_hd__nand3_1 _5227_ (.A(_1170_),
    .B(_1172_),
    .C(_1226_),
    .Y(_1228_));
 sky130_fd_sc_hd__a2bb2o_1 _5228_ (.A1_N(net203),
    .A2_N(_0899_),
    .B1(_1227_),
    .B2(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__a21o_1 _5229_ (.A1(_1166_),
    .A2(_1176_),
    .B1(_1175_),
    .X(_1230_));
 sky130_fd_sc_hd__nand2_1 _5230_ (.A(_1229_),
    .B(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__xor2_1 _5231_ (.A(_1229_),
    .B(_1230_),
    .X(_1232_));
 sky130_fd_sc_hd__and2_1 _5232_ (.A(_1179_),
    .B(_1232_),
    .X(_1233_));
 sky130_fd_sc_hd__xor2_1 _5233_ (.A(_1179_),
    .B(_1232_),
    .X(_1234_));
 sky130_fd_sc_hd__and2_1 _5234_ (.A(_1220_),
    .B(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__nor2_1 _5235_ (.A(_1220_),
    .B(_1234_),
    .Y(_1236_));
 sky130_fd_sc_hd__nor2_2 _5236_ (.A(_1235_),
    .B(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__o21a_2 _5237_ (.A1(_1165_),
    .A2(_1184_),
    .B1(_1183_),
    .X(_1238_));
 sky130_fd_sc_hd__and2b_1 _5238_ (.A_N(_1238_),
    .B(_1237_),
    .X(_1239_));
 sky130_fd_sc_hd__xnor2_4 _5239_ (.A(_1237_),
    .B(_1238_),
    .Y(_1240_));
 sky130_fd_sc_hd__xor2_4 _5240_ (.A(_1203_),
    .B(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__a21o_1 _5241_ (.A1(_1142_),
    .A2(_1188_),
    .B1(_1187_),
    .X(_1242_));
 sky130_fd_sc_hd__xor2_2 _5242_ (.A(_1241_),
    .B(_1242_),
    .X(_1243_));
 sky130_fd_sc_hd__xnor2_1 _5243_ (.A(_1140_),
    .B(_1243_),
    .Y(_1244_));
 sky130_fd_sc_hd__a21oi_1 _5244_ (.A1(_1074_),
    .A2(_1192_),
    .B1(_1191_),
    .Y(_1245_));
 sky130_fd_sc_hd__and2b_1 _5245_ (.A_N(_1245_),
    .B(_1244_),
    .X(_1246_));
 sky130_fd_sc_hd__and2b_1 _5246_ (.A_N(_1244_),
    .B(_1245_),
    .X(_1247_));
 sky130_fd_sc_hd__nor2_2 _5247_ (.A(_1246_),
    .B(_1247_),
    .Y(_1248_));
 sky130_fd_sc_hd__xor2_1 _5248_ (.A(_1244_),
    .B(_1245_),
    .X(_1249_));
 sky130_fd_sc_hd__and4bb_1 _5249_ (.A_N(_1129_),
    .B_N(_1196_),
    .C(_1131_),
    .D(_1195_),
    .X(_1250_));
 sky130_fd_sc_hd__or4_1 _5250_ (.A(_1070_),
    .B(_1129_),
    .C(_1130_),
    .D(_1197_),
    .X(_1251_));
 sky130_fd_sc_hd__a21o_1 _5251_ (.A1(_1128_),
    .A2(_1195_),
    .B1(_1196_),
    .X(_1252_));
 sky130_fd_sc_hd__nand2_1 _5252_ (.A(_1251_),
    .B(_1252_),
    .Y(_1253_));
 sky130_fd_sc_hd__a21o_2 _5253_ (.A1(_1000_),
    .A2(_1250_),
    .B1(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__xnor2_4 _5254_ (.A(_1248_),
    .B(_1254_),
    .Y(_1255_));
 sky130_fd_sc_hd__nor2_1 _5255_ (.A(_1135_),
    .B(_1199_),
    .Y(_1256_));
 sky130_fd_sc_hd__nor2_1 _5256_ (.A(_3620_),
    .B(_1256_),
    .Y(_1257_));
 sky130_fd_sc_hd__xnor2_1 _5257_ (.A(_1255_),
    .B(_1257_),
    .Y(\mul_wb.reg_p[20] ));
 sky130_fd_sc_hd__a21bo_1 _5258_ (.A1(_1205_),
    .A2(_1208_),
    .B1_N(_1206_),
    .X(_1258_));
 sky130_fd_sc_hd__nand2b_1 _5259_ (.A_N(_1219_),
    .B(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__xor2_1 _5260_ (.A(_1219_),
    .B(_1258_),
    .X(_1260_));
 sky130_fd_sc_hd__o21ai_2 _5261_ (.A1(net199),
    .A2(_0862_),
    .B1(_1260_),
    .Y(_1261_));
 sky130_fd_sc_hd__or2_1 _5262_ (.A(_0391_),
    .B(net216),
    .X(_1262_));
 sky130_fd_sc_hd__o211a_1 _5263_ (.A1(_0341_),
    .A2(_0345_),
    .B1(_0821_),
    .C1(_3415_),
    .X(_1263_));
 sky130_fd_sc_hd__nor2_1 _5264_ (.A(net222),
    .B(net220),
    .Y(_1264_));
 sky130_fd_sc_hd__nand2_1 _5265_ (.A(_1263_),
    .B(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__xnor2_2 _5266_ (.A(_1263_),
    .B(_1264_),
    .Y(_1266_));
 sky130_fd_sc_hd__xnor2_1 _5267_ (.A(_1262_),
    .B(_1266_),
    .Y(_1267_));
 sky130_fd_sc_hd__o21ai_2 _5268_ (.A1(_1221_),
    .A2(_1225_),
    .B1(_1224_),
    .Y(_1268_));
 sky130_fd_sc_hd__nand2b_1 _5269_ (.A_N(_1267_),
    .B(_1268_),
    .Y(_1269_));
 sky130_fd_sc_hd__xor2_1 _5270_ (.A(_1267_),
    .B(_1268_),
    .X(_1270_));
 sky130_fd_sc_hd__or2_1 _5271_ (.A(_1227_),
    .B(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__nand2_1 _5272_ (.A(_1227_),
    .B(_1270_),
    .Y(_1272_));
 sky130_fd_sc_hd__nand2_1 _5273_ (.A(_1271_),
    .B(_1272_),
    .Y(_1273_));
 sky130_fd_sc_hd__nor2_1 _5274_ (.A(_1231_),
    .B(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hd__xor2_2 _5275_ (.A(_1231_),
    .B(_1273_),
    .X(_1275_));
 sky130_fd_sc_hd__or2_1 _5276_ (.A(net191),
    .B(net227),
    .X(_1276_));
 sky130_fd_sc_hd__o22a_1 _5277_ (.A1(net197),
    .A2(net237),
    .B1(_0899_),
    .B2(net201),
    .X(_1277_));
 sky130_fd_sc_hd__nor2_1 _5278_ (.A(_1276_),
    .B(_1277_),
    .Y(_1278_));
 sky130_fd_sc_hd__xnor2_2 _5279_ (.A(_1276_),
    .B(_1277_),
    .Y(_1279_));
 sky130_fd_sc_hd__a21boi_2 _5280_ (.A1(_1210_),
    .A2(_1213_),
    .B1_N(_1211_),
    .Y(_1280_));
 sky130_fd_sc_hd__xnor2_2 _5281_ (.A(_1279_),
    .B(_1280_),
    .Y(_1281_));
 sky130_fd_sc_hd__o22a_1 _5282_ (.A1(net189),
    .A2(net221),
    .B1(net218),
    .B2(net224),
    .X(_1282_));
 sky130_fd_sc_hd__nor4_2 _5283_ (.A(net224),
    .B(net189),
    .C(net221),
    .D(net218),
    .Y(_1283_));
 sky130_fd_sc_hd__or2_1 _5284_ (.A(_1282_),
    .B(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__nor2_1 _5285_ (.A(net193),
    .B(net217),
    .Y(_1285_));
 sky130_fd_sc_hd__and2b_1 _5286_ (.A_N(_1284_),
    .B(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__xnor2_2 _5287_ (.A(_1284_),
    .B(_1285_),
    .Y(_1287_));
 sky130_fd_sc_hd__nand2b_1 _5288_ (.A_N(_1281_),
    .B(_1287_),
    .Y(_1288_));
 sky130_fd_sc_hd__xor2_2 _5289_ (.A(_1281_),
    .B(_1287_),
    .X(_1289_));
 sky130_fd_sc_hd__a21bo_1 _5290_ (.A1(_1209_),
    .A2(_1217_),
    .B1_N(_1216_),
    .X(_1290_));
 sky130_fd_sc_hd__and2b_1 _5291_ (.A_N(_1289_),
    .B(_1290_),
    .X(_1291_));
 sky130_fd_sc_hd__xnor2_2 _5292_ (.A(_1289_),
    .B(_1290_),
    .Y(_1292_));
 sky130_fd_sc_hd__xnor2_1 _5293_ (.A(_1275_),
    .B(_1292_),
    .Y(_1293_));
 sky130_fd_sc_hd__o21ba_1 _5294_ (.A1(_1233_),
    .A2(_1235_),
    .B1_N(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__or3b_1 _5295_ (.A(_1233_),
    .B(_1235_),
    .C_N(_1293_),
    .X(_1295_));
 sky130_fd_sc_hd__nand2b_1 _5296_ (.A_N(_1294_),
    .B(_1295_),
    .Y(_1296_));
 sky130_fd_sc_hd__xnor2_2 _5297_ (.A(_1261_),
    .B(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__a21oi_2 _5298_ (.A1(_1203_),
    .A2(_1240_),
    .B1(_1239_),
    .Y(_1298_));
 sky130_fd_sc_hd__and2b_1 _5299_ (.A_N(_1298_),
    .B(_1297_),
    .X(_1299_));
 sky130_fd_sc_hd__xnor2_2 _5300_ (.A(_1297_),
    .B(_1298_),
    .Y(_1300_));
 sky130_fd_sc_hd__xnor2_2 _5301_ (.A(_1201_),
    .B(_1300_),
    .Y(_1301_));
 sky130_fd_sc_hd__a32oi_4 _5302_ (.A1(_1138_),
    .A2(_1139_),
    .A3(_1243_),
    .B1(_1242_),
    .B2(_1241_),
    .Y(_1302_));
 sky130_fd_sc_hd__nor2_1 _5303_ (.A(_1301_),
    .B(_1302_),
    .Y(_1303_));
 sky130_fd_sc_hd__nand2_1 _5304_ (.A(_1301_),
    .B(_1302_),
    .Y(_1304_));
 sky130_fd_sc_hd__xnor2_1 _5305_ (.A(_1301_),
    .B(_1302_),
    .Y(_1305_));
 sky130_fd_sc_hd__inv_2 _5306_ (.A(_1305_),
    .Y(_1306_));
 sky130_fd_sc_hd__a21oi_2 _5307_ (.A1(_1248_),
    .A2(_1254_),
    .B1(_1246_),
    .Y(_1307_));
 sky130_fd_sc_hd__xnor2_4 _5308_ (.A(_1306_),
    .B(_1307_),
    .Y(_1308_));
 sky130_fd_sc_hd__a21o_1 _5309_ (.A1(_1255_),
    .A2(_1256_),
    .B1(_3620_),
    .X(_1309_));
 sky130_fd_sc_hd__xnor2_1 _5310_ (.A(_1308_),
    .B(_1309_),
    .Y(\mul_wb.reg_p[21] ));
 sky130_fd_sc_hd__o22a_1 _5311_ (.A1(net191),
    .A2(net216),
    .B1(_0899_),
    .B2(net197),
    .X(_1310_));
 sky130_fd_sc_hd__and2b_1 _5312_ (.A_N(_1310_),
    .B(_1278_),
    .X(_1311_));
 sky130_fd_sc_hd__xnor2_1 _5313_ (.A(_1278_),
    .B(_1310_),
    .Y(_1312_));
 sky130_fd_sc_hd__o22ai_1 _5314_ (.A1(net222),
    .A2(net218),
    .B1(net227),
    .B2(net189),
    .Y(_1313_));
 sky130_fd_sc_hd__or4_1 _5315_ (.A(net189),
    .B(net222),
    .C(net218),
    .D(net227),
    .X(_1314_));
 sky130_fd_sc_hd__nand2_1 _5316_ (.A(_1313_),
    .B(_1314_),
    .Y(_1315_));
 sky130_fd_sc_hd__nor2_1 _5317_ (.A(net224),
    .B(net217),
    .Y(_1316_));
 sky130_fd_sc_hd__xnor2_1 _5318_ (.A(_1315_),
    .B(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__and2_1 _5319_ (.A(_1312_),
    .B(_1317_),
    .X(_1318_));
 sky130_fd_sc_hd__nor2_1 _5320_ (.A(_1312_),
    .B(_1317_),
    .Y(_1319_));
 sky130_fd_sc_hd__or2_1 _5321_ (.A(_1318_),
    .B(_1319_),
    .X(_1320_));
 sky130_fd_sc_hd__o21a_1 _5322_ (.A1(_1279_),
    .A2(_1280_),
    .B1(_1288_),
    .X(_1321_));
 sky130_fd_sc_hd__or2_1 _5323_ (.A(_1320_),
    .B(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__xnor2_2 _5324_ (.A(_1320_),
    .B(_1321_),
    .Y(_1323_));
 sky130_fd_sc_hd__nor2_1 _5325_ (.A(_0391_),
    .B(net237),
    .Y(_1324_));
 sky130_fd_sc_hd__nand2_1 _5326_ (.A(_0597_),
    .B(_0606_),
    .Y(_1325_));
 sky130_fd_sc_hd__o21ai_1 _5327_ (.A1(net192),
    .A2(_0822_),
    .B1(_1325_),
    .Y(_1326_));
 sky130_fd_sc_hd__or3_1 _5328_ (.A(net193),
    .B(_0822_),
    .C(_1325_),
    .X(_1327_));
 sky130_fd_sc_hd__and2_1 _5329_ (.A(_1326_),
    .B(_1327_),
    .X(_1328_));
 sky130_fd_sc_hd__xnor2_2 _5330_ (.A(_1324_),
    .B(_1328_),
    .Y(_1329_));
 sky130_fd_sc_hd__o21ai_2 _5331_ (.A1(_1262_),
    .A2(_1266_),
    .B1(_1265_),
    .Y(_1330_));
 sky130_fd_sc_hd__and2b_1 _5332_ (.A_N(_1329_),
    .B(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__xor2_2 _5333_ (.A(_1329_),
    .B(_1330_),
    .X(_1332_));
 sky130_fd_sc_hd__nand2_1 _5334_ (.A(_1269_),
    .B(_1271_),
    .Y(_1333_));
 sky130_fd_sc_hd__xor2_2 _5335_ (.A(_1332_),
    .B(_1333_),
    .X(_1334_));
 sky130_fd_sc_hd__xor2_2 _5336_ (.A(_1323_),
    .B(_1334_),
    .X(_1335_));
 sky130_fd_sc_hd__a21oi_2 _5337_ (.A1(_1275_),
    .A2(_1292_),
    .B1(_1274_),
    .Y(_1336_));
 sky130_fd_sc_hd__and2b_1 _5338_ (.A_N(_1336_),
    .B(_1335_),
    .X(_1337_));
 sky130_fd_sc_hd__xnor2_2 _5339_ (.A(_1335_),
    .B(_1336_),
    .Y(_1338_));
 sky130_fd_sc_hd__o21ai_4 _5340_ (.A1(_1283_),
    .A2(_1286_),
    .B1(_1291_),
    .Y(_1339_));
 sky130_fd_sc_hd__or3_1 _5341_ (.A(_1283_),
    .B(_1286_),
    .C(_1291_),
    .X(_1340_));
 sky130_fd_sc_hd__o2bb2a_1 _5342_ (.A1_N(_1339_),
    .A2_N(_1340_),
    .B1(_0346_),
    .B2(_0862_),
    .X(_1341_));
 sky130_fd_sc_hd__inv_2 _5343_ (.A(_1341_),
    .Y(_1342_));
 sky130_fd_sc_hd__xnor2_1 _5344_ (.A(_1338_),
    .B(_1341_),
    .Y(_1343_));
 sky130_fd_sc_hd__a21oi_1 _5345_ (.A1(_1261_),
    .A2(_1295_),
    .B1(_1294_),
    .Y(_1344_));
 sky130_fd_sc_hd__nand2b_1 _5346_ (.A_N(_1344_),
    .B(_1343_),
    .Y(_1345_));
 sky130_fd_sc_hd__xor2_1 _5347_ (.A(_1343_),
    .B(_1344_),
    .X(_1346_));
 sky130_fd_sc_hd__or2_1 _5348_ (.A(_1259_),
    .B(_1346_),
    .X(_1347_));
 sky130_fd_sc_hd__nand2_1 _5349_ (.A(_1259_),
    .B(_1346_),
    .Y(_1348_));
 sky130_fd_sc_hd__and2_2 _5350_ (.A(_1347_),
    .B(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__a21oi_2 _5351_ (.A1(_1201_),
    .A2(_1300_),
    .B1(_1299_),
    .Y(_1350_));
 sky130_fd_sc_hd__and2b_1 _5352_ (.A_N(_1350_),
    .B(_1349_),
    .X(_1351_));
 sky130_fd_sc_hd__xnor2_4 _5353_ (.A(_1349_),
    .B(_1350_),
    .Y(_1352_));
 sky130_fd_sc_hd__o21a_1 _5354_ (.A1(_1246_),
    .A2(_1303_),
    .B1(_1304_),
    .X(_1353_));
 sky130_fd_sc_hd__a31o_2 _5355_ (.A1(_1248_),
    .A2(_1254_),
    .A3(_1306_),
    .B1(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__xor2_4 _5356_ (.A(_1352_),
    .B(_1354_),
    .X(_1355_));
 sky130_fd_sc_hd__or4b_2 _5357_ (.A(_1135_),
    .B(_1199_),
    .C(_1308_),
    .D_N(_1255_),
    .X(_1356_));
 sky130_fd_sc_hd__nand2_1 _5358_ (.A(net252),
    .B(_1356_),
    .Y(_1357_));
 sky130_fd_sc_hd__xnor2_1 _5359_ (.A(_1355_),
    .B(_1357_),
    .Y(\mul_wb.reg_p[22] ));
 sky130_fd_sc_hd__o21a_1 _5360_ (.A1(_1355_),
    .A2(_1356_),
    .B1(net252),
    .X(_1358_));
 sky130_fd_sc_hd__o22ai_1 _5361_ (.A1(_0598_),
    .A2(net218),
    .B1(net216),
    .B2(net189),
    .Y(_1359_));
 sky130_fd_sc_hd__or4_1 _5362_ (.A(net189),
    .B(net221),
    .C(net218),
    .D(net216),
    .X(_1360_));
 sky130_fd_sc_hd__nand2_1 _5363_ (.A(_1359_),
    .B(_1360_),
    .Y(_1361_));
 sky130_fd_sc_hd__nor2_1 _5364_ (.A(_0535_),
    .B(net217),
    .Y(_1362_));
 sky130_fd_sc_hd__xor2_1 _5365_ (.A(_1361_),
    .B(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__or3_1 _5366_ (.A(_0442_),
    .B(net237),
    .C(_1363_),
    .X(_1364_));
 sky130_fd_sc_hd__o21ai_1 _5367_ (.A1(_0442_),
    .A2(net237),
    .B1(_1363_),
    .Y(_1365_));
 sky130_fd_sc_hd__and2_1 _5368_ (.A(_1364_),
    .B(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__o21ai_2 _5369_ (.A1(_1311_),
    .A2(_1318_),
    .B1(_1366_),
    .Y(_1367_));
 sky130_fd_sc_hd__or3_1 _5370_ (.A(_1311_),
    .B(_1318_),
    .C(_1366_),
    .X(_1368_));
 sky130_fd_sc_hd__nand2_2 _5371_ (.A(_1367_),
    .B(_1368_),
    .Y(_1369_));
 sky130_fd_sc_hd__a21bo_1 _5372_ (.A1(_1324_),
    .A2(_1328_),
    .B1_N(_1327_),
    .X(_1370_));
 sky130_fd_sc_hd__o22ai_1 _5373_ (.A1(net220),
    .A2(net227),
    .B1(_0822_),
    .B2(net223),
    .Y(_1371_));
 sky130_fd_sc_hd__or4_1 _5374_ (.A(net224),
    .B(net220),
    .C(net227),
    .D(_0822_),
    .X(_1372_));
 sky130_fd_sc_hd__a2bb2o_1 _5375_ (.A1_N(_0391_),
    .A2_N(_0899_),
    .B1(_1371_),
    .B2(_1372_),
    .X(_1373_));
 sky130_fd_sc_hd__nand2_1 _5376_ (.A(_1370_),
    .B(_1373_),
    .Y(_1374_));
 sky130_fd_sc_hd__xnor2_2 _5377_ (.A(_1370_),
    .B(_1373_),
    .Y(_1375_));
 sky130_fd_sc_hd__inv_2 _5378_ (.A(_1375_),
    .Y(_1376_));
 sky130_fd_sc_hd__nor2_1 _5379_ (.A(_1269_),
    .B(_1332_),
    .Y(_1377_));
 sky130_fd_sc_hd__nor2_1 _5380_ (.A(_1331_),
    .B(_1377_),
    .Y(_1378_));
 sky130_fd_sc_hd__xnor2_2 _5381_ (.A(_1375_),
    .B(_1378_),
    .Y(_1379_));
 sky130_fd_sc_hd__xnor2_4 _5382_ (.A(_1369_),
    .B(_1379_),
    .Y(_1380_));
 sky130_fd_sc_hd__o22a_2 _5383_ (.A1(_1271_),
    .A2(_1332_),
    .B1(_1334_),
    .B2(_1323_),
    .X(_1381_));
 sky130_fd_sc_hd__or2_1 _5384_ (.A(_1380_),
    .B(_1381_),
    .X(_1382_));
 sky130_fd_sc_hd__xnor2_4 _5385_ (.A(_1380_),
    .B(_1381_),
    .Y(_1383_));
 sky130_fd_sc_hd__a21bo_1 _5386_ (.A1(_1313_),
    .A2(_1316_),
    .B1_N(_1314_),
    .X(_1384_));
 sky130_fd_sc_hd__and2b_1 _5387_ (.A_N(_1322_),
    .B(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__xor2_1 _5388_ (.A(_1322_),
    .B(_1384_),
    .X(_1386_));
 sky130_fd_sc_hd__o21a_2 _5389_ (.A1(net193),
    .A2(_0862_),
    .B1(_1386_),
    .X(_1387_));
 sky130_fd_sc_hd__xnor2_4 _5390_ (.A(_1383_),
    .B(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__a21oi_4 _5391_ (.A1(_1338_),
    .A2(_1342_),
    .B1(_1337_),
    .Y(_1389_));
 sky130_fd_sc_hd__xnor2_4 _5392_ (.A(_1388_),
    .B(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__or2_1 _5393_ (.A(_1339_),
    .B(_1390_),
    .X(_1391_));
 sky130_fd_sc_hd__xnor2_4 _5394_ (.A(_1339_),
    .B(_1390_),
    .Y(_1392_));
 sky130_fd_sc_hd__nand2_2 _5395_ (.A(_1345_),
    .B(_1347_),
    .Y(_1393_));
 sky130_fd_sc_hd__nand2b_1 _5396_ (.A_N(_1393_),
    .B(_1392_),
    .Y(_1394_));
 sky130_fd_sc_hd__and2b_1 _5397_ (.A_N(_1392_),
    .B(_1393_),
    .X(_1395_));
 sky130_fd_sc_hd__xor2_4 _5398_ (.A(_1392_),
    .B(_1393_),
    .X(_1396_));
 sky130_fd_sc_hd__inv_2 _5399_ (.A(_1396_),
    .Y(_1397_));
 sky130_fd_sc_hd__a21oi_2 _5400_ (.A1(_1352_),
    .A2(_1354_),
    .B1(_1351_),
    .Y(_1398_));
 sky130_fd_sc_hd__xnor2_4 _5401_ (.A(_1396_),
    .B(_1398_),
    .Y(_1399_));
 sky130_fd_sc_hd__xnor2_1 _5402_ (.A(_1358_),
    .B(_1399_),
    .Y(\mul_wb.reg_p[23] ));
 sky130_fd_sc_hd__o22a_1 _5403_ (.A1(net218),
    .A2(net227),
    .B1(net237),
    .B2(net189),
    .X(_1400_));
 sky130_fd_sc_hd__or4_1 _5404_ (.A(net189),
    .B(net218),
    .C(net227),
    .D(net237),
    .X(_1401_));
 sky130_fd_sc_hd__and2b_1 _5405_ (.A_N(_1400_),
    .B(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__nor2_1 _5406_ (.A(net221),
    .B(net217),
    .Y(_1403_));
 sky130_fd_sc_hd__xnor2_1 _5407_ (.A(_1402_),
    .B(_1403_),
    .Y(_1404_));
 sky130_fd_sc_hd__o21a_1 _5408_ (.A1(_0442_),
    .A2(_0899_),
    .B1(_1404_),
    .X(_1405_));
 sky130_fd_sc_hd__or2_1 _5409_ (.A(_1364_),
    .B(_1405_),
    .X(_1406_));
 sky130_fd_sc_hd__nand2_1 _5410_ (.A(_1364_),
    .B(_1405_),
    .Y(_1407_));
 sky130_fd_sc_hd__nand2_1 _5411_ (.A(_1406_),
    .B(_1407_),
    .Y(_1408_));
 sky130_fd_sc_hd__nand2_1 _5412_ (.A(_1331_),
    .B(_1376_),
    .Y(_1409_));
 sky130_fd_sc_hd__a22o_1 _5413_ (.A1(_0606_),
    .A2(_0752_),
    .B1(_0821_),
    .B2(_0536_),
    .X(_1410_));
 sky130_fd_sc_hd__or4_1 _5414_ (.A(_0535_),
    .B(_0607_),
    .C(net216),
    .D(_0822_),
    .X(_1411_));
 sky130_fd_sc_hd__nand2_1 _5415_ (.A(_1410_),
    .B(_1411_),
    .Y(_1412_));
 sky130_fd_sc_hd__or2_1 _5416_ (.A(_1372_),
    .B(_1412_),
    .X(_1413_));
 sky130_fd_sc_hd__nand2_1 _5417_ (.A(_1372_),
    .B(_1412_),
    .Y(_1414_));
 sky130_fd_sc_hd__nand2_1 _5418_ (.A(_1413_),
    .B(_1414_),
    .Y(_1415_));
 sky130_fd_sc_hd__nor2_1 _5419_ (.A(_1409_),
    .B(_1415_),
    .Y(_1416_));
 sky130_fd_sc_hd__and3_1 _5420_ (.A(_1374_),
    .B(_1409_),
    .C(_1415_),
    .X(_1417_));
 sky130_fd_sc_hd__or2_1 _5421_ (.A(_1374_),
    .B(_1415_),
    .X(_1418_));
 sky130_fd_sc_hd__or3b_1 _5422_ (.A(_1416_),
    .B(_1417_),
    .C_N(_1418_),
    .X(_1419_));
 sky130_fd_sc_hd__nor2_1 _5423_ (.A(_1408_),
    .B(_1419_),
    .Y(_1420_));
 sky130_fd_sc_hd__xor2_1 _5424_ (.A(_1408_),
    .B(_1419_),
    .X(_1421_));
 sky130_fd_sc_hd__o2bb2a_1 _5425_ (.A1_N(_1376_),
    .A2_N(_1377_),
    .B1(_1379_),
    .B2(_1369_),
    .X(_1422_));
 sky130_fd_sc_hd__and2b_1 _5426_ (.A_N(_1422_),
    .B(_1421_),
    .X(_1423_));
 sky130_fd_sc_hd__xnor2_1 _5427_ (.A(_1421_),
    .B(_1422_),
    .Y(_1424_));
 sky130_fd_sc_hd__a21bo_1 _5428_ (.A1(_1359_),
    .A2(_1362_),
    .B1_N(_1360_),
    .X(_1425_));
 sky130_fd_sc_hd__nand2b_1 _5429_ (.A_N(_1367_),
    .B(_1425_),
    .Y(_1426_));
 sky130_fd_sc_hd__xnor2_1 _5430_ (.A(_1367_),
    .B(_1425_),
    .Y(_1427_));
 sky130_fd_sc_hd__nor2_1 _5431_ (.A(net224),
    .B(_0862_),
    .Y(_1428_));
 sky130_fd_sc_hd__o21a_1 _5432_ (.A1(_1427_),
    .A2(_1428_),
    .B1(_1424_),
    .X(_1429_));
 sky130_fd_sc_hd__nor3_1 _5433_ (.A(_1424_),
    .B(_1427_),
    .C(_1428_),
    .Y(_1430_));
 sky130_fd_sc_hd__nor2_1 _5434_ (.A(_1429_),
    .B(_1430_),
    .Y(_1431_));
 sky130_fd_sc_hd__o21a_1 _5435_ (.A1(_1383_),
    .A2(_1387_),
    .B1(_1382_),
    .X(_1432_));
 sky130_fd_sc_hd__or3_1 _5436_ (.A(_1429_),
    .B(_1430_),
    .C(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__xnor2_1 _5437_ (.A(_1431_),
    .B(_1432_),
    .Y(_1434_));
 sky130_fd_sc_hd__nand2_1 _5438_ (.A(_1385_),
    .B(_1434_),
    .Y(_1435_));
 sky130_fd_sc_hd__or2_1 _5439_ (.A(_1385_),
    .B(_1434_),
    .X(_1436_));
 sky130_fd_sc_hd__and2_1 _5440_ (.A(_1435_),
    .B(_1436_),
    .X(_1437_));
 sky130_fd_sc_hd__o21a_1 _5441_ (.A1(_1388_),
    .A2(_1389_),
    .B1(_1391_),
    .X(_1438_));
 sky130_fd_sc_hd__nand2b_1 _5442_ (.A_N(_1438_),
    .B(_1437_),
    .Y(_1439_));
 sky130_fd_sc_hd__xnor2_1 _5443_ (.A(_1437_),
    .B(_1438_),
    .Y(_1440_));
 sky130_fd_sc_hd__inv_2 _5444_ (.A(_1440_),
    .Y(_1441_));
 sky130_fd_sc_hd__and2_1 _5445_ (.A(_1352_),
    .B(_1397_),
    .X(_1442_));
 sky130_fd_sc_hd__a221oi_4 _5446_ (.A1(_1351_),
    .A2(_1394_),
    .B1(_1442_),
    .B2(_1353_),
    .C1(_1395_),
    .Y(_1443_));
 sky130_fd_sc_hd__or4bb_2 _5447_ (.A(_1249_),
    .B(_1305_),
    .C_N(_1352_),
    .D_N(_1397_),
    .X(_1444_));
 sky130_fd_sc_hd__inv_2 _5448_ (.A(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__a21oi_1 _5449_ (.A1(_1251_),
    .A2(_1252_),
    .B1(_1444_),
    .Y(_1446_));
 sky130_fd_sc_hd__a31oi_4 _5450_ (.A1(_1000_),
    .A2(_1250_),
    .A3(_1445_),
    .B1(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__nand2_1 _5451_ (.A(_1443_),
    .B(_1447_),
    .Y(_1448_));
 sky130_fd_sc_hd__a21o_1 _5452_ (.A1(_1443_),
    .A2(_1447_),
    .B1(_1441_),
    .X(_1449_));
 sky130_fd_sc_hd__xnor2_2 _5453_ (.A(_1441_),
    .B(_1448_),
    .Y(_1450_));
 sky130_fd_sc_hd__or3b_1 _5454_ (.A(_1355_),
    .B(_1356_),
    .C_N(_1399_),
    .X(_1451_));
 sky130_fd_sc_hd__nand2_1 _5455_ (.A(net252),
    .B(_1451_),
    .Y(_1452_));
 sky130_fd_sc_hd__xnor2_1 _5456_ (.A(_1450_),
    .B(_1452_),
    .Y(\mul_wb.reg_p[24] ));
 sky130_fd_sc_hd__a2bb2o_1 _5457_ (.A1_N(_0607_),
    .A2_N(net237),
    .B1(_0821_),
    .B2(_0597_),
    .X(_1453_));
 sky130_fd_sc_hd__or3_2 _5458_ (.A(_3396_),
    .B(_0822_),
    .C(_1325_),
    .X(_1454_));
 sky130_fd_sc_hd__nand2_1 _5459_ (.A(_1453_),
    .B(_1454_),
    .Y(_1455_));
 sky130_fd_sc_hd__nor2_1 _5460_ (.A(_1413_),
    .B(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__and3_1 _5461_ (.A(_1411_),
    .B(_1413_),
    .C(_1455_),
    .X(_1457_));
 sky130_fd_sc_hd__or2_1 _5462_ (.A(_1411_),
    .B(_1455_),
    .X(_1458_));
 sky130_fd_sc_hd__or3b_1 _5463_ (.A(_1456_),
    .B(_1457_),
    .C_N(_1458_),
    .X(_1459_));
 sky130_fd_sc_hd__or2_1 _5464_ (.A(_1418_),
    .B(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__nand2_1 _5465_ (.A(_1418_),
    .B(_1459_),
    .Y(_1461_));
 sky130_fd_sc_hd__nand2_1 _5466_ (.A(_1460_),
    .B(_1461_),
    .Y(_1462_));
 sky130_fd_sc_hd__o22a_1 _5467_ (.A1(net218),
    .A2(net216),
    .B1(_0899_),
    .B2(net189),
    .X(_1463_));
 sky130_fd_sc_hd__or2_1 _5468_ (.A(net227),
    .B(net217),
    .X(_1464_));
 sky130_fd_sc_hd__xnor2_1 _5469_ (.A(_1463_),
    .B(_1464_),
    .Y(_1465_));
 sky130_fd_sc_hd__xor2_1 _5470_ (.A(_1462_),
    .B(_1465_),
    .X(_1466_));
 sky130_fd_sc_hd__o21a_1 _5471_ (.A1(_1416_),
    .A2(_1420_),
    .B1(_1466_),
    .X(_1467_));
 sky130_fd_sc_hd__nor3_1 _5472_ (.A(_1416_),
    .B(_1420_),
    .C(_1466_),
    .Y(_1468_));
 sky130_fd_sc_hd__nor2_1 _5473_ (.A(_1467_),
    .B(_1468_),
    .Y(_1469_));
 sky130_fd_sc_hd__a21bo_1 _5474_ (.A1(_1402_),
    .A2(_1403_),
    .B1_N(_1401_),
    .X(_1470_));
 sky130_fd_sc_hd__or3b_1 _5475_ (.A(_1364_),
    .B(_1405_),
    .C_N(_1470_),
    .X(_1471_));
 sky130_fd_sc_hd__xnor2_1 _5476_ (.A(_1406_),
    .B(_1470_),
    .Y(_1472_));
 sky130_fd_sc_hd__a31o_1 _5477_ (.A1(net269),
    .A2(net242),
    .A3(_0536_),
    .B1(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__xor2_1 _5478_ (.A(_1469_),
    .B(_1473_),
    .X(_1474_));
 sky130_fd_sc_hd__o21ai_1 _5479_ (.A1(_1423_),
    .A2(_1429_),
    .B1(_1474_),
    .Y(_1475_));
 sky130_fd_sc_hd__or3_1 _5480_ (.A(_1423_),
    .B(_1429_),
    .C(_1474_),
    .X(_1476_));
 sky130_fd_sc_hd__and2_1 _5481_ (.A(_1475_),
    .B(_1476_),
    .X(_1477_));
 sky130_fd_sc_hd__nand2b_1 _5482_ (.A_N(_1426_),
    .B(_1477_),
    .Y(_1478_));
 sky130_fd_sc_hd__xor2_1 _5483_ (.A(_1426_),
    .B(_1477_),
    .X(_1479_));
 sky130_fd_sc_hd__nand2_1 _5484_ (.A(_1433_),
    .B(_1435_),
    .Y(_1480_));
 sky130_fd_sc_hd__nand2b_1 _5485_ (.A_N(_1479_),
    .B(_1480_),
    .Y(_1481_));
 sky130_fd_sc_hd__and3_1 _5486_ (.A(_1433_),
    .B(_1435_),
    .C(_1479_),
    .X(_1482_));
 sky130_fd_sc_hd__xnor2_1 _5487_ (.A(_1479_),
    .B(_1480_),
    .Y(_1483_));
 sky130_fd_sc_hd__and3_1 _5488_ (.A(_1439_),
    .B(_1449_),
    .C(_1483_),
    .X(_1484_));
 sky130_fd_sc_hd__a21oi_1 _5489_ (.A1(_1439_),
    .A2(_1449_),
    .B1(_1483_),
    .Y(_1485_));
 sky130_fd_sc_hd__or2_1 _5490_ (.A(_1484_),
    .B(_1485_),
    .X(_1486_));
 sky130_fd_sc_hd__o21ai_1 _5491_ (.A1(_1450_),
    .A2(_1451_),
    .B1(net252),
    .Y(_1487_));
 sky130_fd_sc_hd__xnor2_1 _5492_ (.A(_1486_),
    .B(_1487_),
    .Y(\mul_wb.reg_p[25] ));
 sky130_fd_sc_hd__o22a_1 _5493_ (.A1(net227),
    .A2(_0822_),
    .B1(_0899_),
    .B2(_0607_),
    .X(_1488_));
 sky130_fd_sc_hd__a21oi_1 _5494_ (.A1(_1454_),
    .A2(_1458_),
    .B1(_1488_),
    .Y(_1489_));
 sky130_fd_sc_hd__a31o_1 _5495_ (.A1(_1454_),
    .A2(_1458_),
    .A3(_1488_),
    .B1(_1456_),
    .X(_1490_));
 sky130_fd_sc_hd__or2_1 _5496_ (.A(_1489_),
    .B(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__o22ai_1 _5497_ (.A1(net217),
    .A2(net216),
    .B1(net237),
    .B2(net218),
    .Y(_1492_));
 sky130_fd_sc_hd__or4_1 _5498_ (.A(net218),
    .B(net217),
    .C(net216),
    .D(net237),
    .X(_1493_));
 sky130_fd_sc_hd__nand2_1 _5499_ (.A(_1492_),
    .B(_1493_),
    .Y(_1494_));
 sky130_fd_sc_hd__xnor2_1 _5500_ (.A(_1491_),
    .B(_1494_),
    .Y(_1495_));
 sky130_fd_sc_hd__o21a_1 _5501_ (.A1(_1462_),
    .A2(_1465_),
    .B1(_1460_),
    .X(_1496_));
 sky130_fd_sc_hd__nor2_1 _5502_ (.A(_1495_),
    .B(_1496_),
    .Y(_1497_));
 sky130_fd_sc_hd__xnor2_1 _5503_ (.A(_1495_),
    .B(_1496_),
    .Y(_1498_));
 sky130_fd_sc_hd__o22a_1 _5504_ (.A1(net221),
    .A2(_0862_),
    .B1(_1463_),
    .B2(_1464_),
    .X(_1499_));
 sky130_fd_sc_hd__nor2_1 _5505_ (.A(_1498_),
    .B(_1499_),
    .Y(_1500_));
 sky130_fd_sc_hd__and2_1 _5506_ (.A(_1498_),
    .B(_1499_),
    .X(_1501_));
 sky130_fd_sc_hd__or2_1 _5507_ (.A(_1500_),
    .B(_1501_),
    .X(_1502_));
 sky130_fd_sc_hd__a21oi_1 _5508_ (.A1(_1469_),
    .A2(_1473_),
    .B1(_1467_),
    .Y(_1503_));
 sky130_fd_sc_hd__nor2_1 _5509_ (.A(_1502_),
    .B(_1503_),
    .Y(_1504_));
 sky130_fd_sc_hd__xnor2_1 _5510_ (.A(_1502_),
    .B(_1503_),
    .Y(_1505_));
 sky130_fd_sc_hd__nor2_1 _5511_ (.A(_1471_),
    .B(_1505_),
    .Y(_1506_));
 sky130_fd_sc_hd__and2_1 _5512_ (.A(_1471_),
    .B(_1505_),
    .X(_1507_));
 sky130_fd_sc_hd__or2_1 _5513_ (.A(_1506_),
    .B(_1507_),
    .X(_1508_));
 sky130_fd_sc_hd__a21oi_1 _5514_ (.A1(_1475_),
    .A2(_1478_),
    .B1(_1508_),
    .Y(_1509_));
 sky130_fd_sc_hd__and3_1 _5515_ (.A(_1475_),
    .B(_1478_),
    .C(_1508_),
    .X(_1510_));
 sky130_fd_sc_hd__nor2_1 _5516_ (.A(_1509_),
    .B(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__inv_2 _5517_ (.A(_1511_),
    .Y(_1512_));
 sky130_fd_sc_hd__nand2_1 _5518_ (.A(_1440_),
    .B(_1483_),
    .Y(_1513_));
 sky130_fd_sc_hd__a21o_1 _5519_ (.A1(_1443_),
    .A2(_1447_),
    .B1(_1513_),
    .X(_1514_));
 sky130_fd_sc_hd__a21o_1 _5520_ (.A1(_1439_),
    .A2(_1481_),
    .B1(_1482_),
    .X(_1515_));
 sky130_fd_sc_hd__a21o_1 _5521_ (.A1(_1514_),
    .A2(_1515_),
    .B1(_1512_),
    .X(_1516_));
 sky130_fd_sc_hd__nand3_1 _5522_ (.A(_1512_),
    .B(_1514_),
    .C(_1515_),
    .Y(_1517_));
 sky130_fd_sc_hd__and2_1 _5523_ (.A(_1516_),
    .B(_1517_),
    .X(_1518_));
 sky130_fd_sc_hd__o31a_1 _5524_ (.A1(_1450_),
    .A2(_1451_),
    .A3(_1486_),
    .B1(net698),
    .X(_1519_));
 sky130_fd_sc_hd__xor2_1 _5525_ (.A(_1518_),
    .B(_1519_),
    .X(\mul_wb.reg_p[26] ));
 sky130_fd_sc_hd__nor2_1 _5526_ (.A(_1458_),
    .B(_1488_),
    .Y(_1520_));
 sky130_fd_sc_hd__a2bb2o_1 _5527_ (.A1_N(_1454_),
    .A2_N(_1488_),
    .B1(_0752_),
    .B2(_0821_),
    .X(_1521_));
 sky130_fd_sc_hd__or4_1 _5528_ (.A(net216),
    .B(_0822_),
    .C(_1454_),
    .D(_1488_),
    .X(_1522_));
 sky130_fd_sc_hd__nand2_1 _5529_ (.A(_1521_),
    .B(_1522_),
    .Y(_1523_));
 sky130_fd_sc_hd__nor2_1 _5530_ (.A(_1520_),
    .B(_1523_),
    .Y(_1524_));
 sky130_fd_sc_hd__o22a_1 _5531_ (.A1(net217),
    .A2(net237),
    .B1(_0899_),
    .B2(net218),
    .X(_1525_));
 sky130_fd_sc_hd__xnor2_1 _5532_ (.A(_1524_),
    .B(_1525_),
    .Y(_1526_));
 sky130_fd_sc_hd__o21ba_1 _5533_ (.A1(_1491_),
    .A2(_1494_),
    .B1_N(_1456_),
    .X(_1527_));
 sky130_fd_sc_hd__and2b_1 _5534_ (.A_N(_1527_),
    .B(_1526_),
    .X(_1528_));
 sky130_fd_sc_hd__xnor2_1 _5535_ (.A(_1526_),
    .B(_1527_),
    .Y(_1529_));
 sky130_fd_sc_hd__o21ai_1 _5536_ (.A1(net227),
    .A2(_0862_),
    .B1(_1493_),
    .Y(_1530_));
 sky130_fd_sc_hd__xor2_1 _5537_ (.A(_1529_),
    .B(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__o21ai_1 _5538_ (.A1(_1497_),
    .A2(_1500_),
    .B1(_1531_),
    .Y(_1532_));
 sky130_fd_sc_hd__or3_1 _5539_ (.A(_1497_),
    .B(_1500_),
    .C(_1531_),
    .X(_1533_));
 sky130_fd_sc_hd__and2_1 _5540_ (.A(_1532_),
    .B(_1533_),
    .X(_1534_));
 sky130_fd_sc_hd__or3_1 _5541_ (.A(_1504_),
    .B(_1506_),
    .C(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__o21ai_1 _5542_ (.A1(_1504_),
    .A2(_1506_),
    .B1(_1534_),
    .Y(_1536_));
 sky130_fd_sc_hd__nand2_2 _5543_ (.A(_1535_),
    .B(_1536_),
    .Y(_1537_));
 sky130_fd_sc_hd__and2b_1 _5544_ (.A_N(_1509_),
    .B(_1516_),
    .X(_1538_));
 sky130_fd_sc_hd__xnor2_2 _5545_ (.A(_1537_),
    .B(_1538_),
    .Y(_1539_));
 sky130_fd_sc_hd__a2111oi_1 _5546_ (.A1(_1516_),
    .A2(_1517_),
    .B1(_1450_),
    .C1(_1484_),
    .D1(_1485_),
    .Y(_1540_));
 sky130_fd_sc_hd__and4bb_1 _5547_ (.A_N(_1355_),
    .B_N(_1356_),
    .C(_1399_),
    .D(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__nor2_1 _5548_ (.A(_3620_),
    .B(_1541_),
    .Y(_1542_));
 sky130_fd_sc_hd__xnor2_1 _5549_ (.A(_1539_),
    .B(_1542_),
    .Y(\mul_wb.reg_p[27] ));
 sky130_fd_sc_hd__nor2_1 _5550_ (.A(net217),
    .B(_0899_),
    .Y(_1543_));
 sky130_fd_sc_hd__a31o_1 _5551_ (.A1(net249),
    .A2(_0821_),
    .A3(_1522_),
    .B1(_1543_),
    .X(_1544_));
 sky130_fd_sc_hd__o21bai_1 _5552_ (.A1(_1523_),
    .A2(_1525_),
    .B1_N(_1520_),
    .Y(_1545_));
 sky130_fd_sc_hd__xor2_1 _5553_ (.A(_1544_),
    .B(_1545_),
    .X(_1546_));
 sky130_fd_sc_hd__o21ba_1 _5554_ (.A1(net216),
    .A2(_0862_),
    .B1_N(_1546_),
    .X(_1547_));
 sky130_fd_sc_hd__a21oi_1 _5555_ (.A1(_1529_),
    .A2(_1530_),
    .B1(_1528_),
    .Y(_1548_));
 sky130_fd_sc_hd__xnor2_1 _5556_ (.A(_1547_),
    .B(_1548_),
    .Y(_1549_));
 sky130_fd_sc_hd__nor2_1 _5557_ (.A(_1532_),
    .B(_1549_),
    .Y(_1550_));
 sky130_fd_sc_hd__and2_1 _5558_ (.A(_1532_),
    .B(_1549_),
    .X(_1551_));
 sky130_fd_sc_hd__or2_1 _5559_ (.A(_1550_),
    .B(_1551_),
    .X(_1552_));
 sky130_fd_sc_hd__a21boi_1 _5560_ (.A1(_1509_),
    .A2(_1535_),
    .B1_N(_1536_),
    .Y(_1553_));
 sky130_fd_sc_hd__or3_1 _5561_ (.A(_1512_),
    .B(_1514_),
    .C(_1537_),
    .X(_1554_));
 sky130_fd_sc_hd__o311a_1 _5562_ (.A1(_1512_),
    .A2(_1515_),
    .A3(_1537_),
    .B1(_1553_),
    .C1(_1554_),
    .X(_1555_));
 sky130_fd_sc_hd__nor2_1 _5563_ (.A(_1552_),
    .B(_1555_),
    .Y(_1556_));
 sky130_fd_sc_hd__xnor2_1 _5564_ (.A(_1552_),
    .B(_1555_),
    .Y(_1557_));
 sky130_fd_sc_hd__a21oi_1 _5565_ (.A1(_1539_),
    .A2(_1541_),
    .B1(_3620_),
    .Y(_1558_));
 sky130_fd_sc_hd__xnor2_1 _5566_ (.A(_1557_),
    .B(_1558_),
    .Y(\mul_wb.reg_p[28] ));
 sky130_fd_sc_hd__o221a_1 _5567_ (.A1(_3396_),
    .A2(_0862_),
    .B1(_0899_),
    .B2(net244),
    .C1(_1522_),
    .X(_1559_));
 sky130_fd_sc_hd__a21boi_1 _5568_ (.A1(_1544_),
    .A2(_1545_),
    .B1_N(_1559_),
    .Y(_1560_));
 sky130_fd_sc_hd__o21ai_1 _5569_ (.A1(_1547_),
    .A2(_1548_),
    .B1(_1560_),
    .Y(_1561_));
 sky130_fd_sc_hd__or3_1 _5570_ (.A(_1550_),
    .B(_1556_),
    .C(_1561_),
    .X(_1562_));
 sky130_fd_sc_hd__a31o_1 _5571_ (.A1(_1539_),
    .A2(_1541_),
    .A3(_1557_),
    .B1(_3620_),
    .X(_1563_));
 sky130_fd_sc_hd__xnor2_1 _5572_ (.A(_1562_),
    .B(_1563_),
    .Y(\mul_wb.reg_p[29] ));
 sky130_fd_sc_hd__and4bb_1 _5573_ (.A_N(_1550_),
    .B_N(_1561_),
    .C(_1552_),
    .D(_1555_),
    .X(_1564_));
 sky130_fd_sc_hd__a31oi_2 _5574_ (.A1(_1539_),
    .A2(_1541_),
    .A3(_1564_),
    .B1(_3620_),
    .Y(\mul_wb.reg_p[31] ));
 sky130_fd_sc_hd__a31o_1 _5575_ (.A1(net269),
    .A2(_3397_),
    .A3(net970),
    .B1(\mul_wb.reg_p[31] ),
    .X(\mul_wb.reg_p[30] ));
 sky130_fd_sc_hd__or4_4 _5576_ (.A(\mul_la.reg_b0[1] ),
    .B(\mul_la.lob_4.B[0] ),
    .C(\mul_la.reg_b0[2] ),
    .D(\mul_la.reg_b0[3] ),
    .X(_1565_));
 sky130_fd_sc_hd__or2_4 _5577_ (.A(\mul_la.reg_b0[4] ),
    .B(\mul_la.reg_b0[5] ),
    .X(_1566_));
 sky130_fd_sc_hd__or2_2 _5578_ (.A(\mul_la.reg_b0[6] ),
    .B(\mul_la.reg_b0[7] ),
    .X(_1567_));
 sky130_fd_sc_hd__or2_1 _5579_ (.A(\mul_la.reg_b0[8] ),
    .B(\mul_la.reg_b0[9] ),
    .X(_1568_));
 sky130_fd_sc_hd__or4_1 _5580_ (.A(\mul_la.reg_b0[8] ),
    .B(\mul_la.reg_b0[9] ),
    .C(\mul_la.reg_b0[10] ),
    .D(\mul_la.reg_b0[11] ),
    .X(_1569_));
 sky130_fd_sc_hd__nor4_2 _5581_ (.A(_1565_),
    .B(_1566_),
    .C(_1567_),
    .D(_1569_),
    .Y(_1570_));
 sky130_fd_sc_hd__nor2_2 _5582_ (.A(\mul_la.reg_b0[12] ),
    .B(\mul_la.reg_b0[13] ),
    .Y(_1571_));
 sky130_fd_sc_hd__and2_1 _5583_ (.A(_1570_),
    .B(_1571_),
    .X(_1572_));
 sky130_fd_sc_hd__a21boi_4 _5584_ (.A1(_1570_),
    .A2(_1571_),
    .B1_N(net254),
    .Y(_1573_));
 sky130_fd_sc_hd__and2_1 _5585_ (.A(net254),
    .B(_3376_),
    .X(_1574_));
 sky130_fd_sc_hd__nand2_2 _5586_ (.A(\mul_la.reg_b0[15] ),
    .B(_3376_),
    .Y(_1575_));
 sky130_fd_sc_hd__a21o_1 _5587_ (.A1(_1570_),
    .A2(_1571_),
    .B1(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__o21ai_4 _5588_ (.A1(_3376_),
    .A2(_1573_),
    .B1(_1576_),
    .Y(_1577_));
 sky130_fd_sc_hd__o41a_4 _5589_ (.A1(_1565_),
    .A2(_1566_),
    .A3(_1567_),
    .A4(_1569_),
    .B1(net254),
    .X(_1578_));
 sky130_fd_sc_hd__and2_1 _5590_ (.A(net254),
    .B(\mul_la.reg_b0[12] ),
    .X(_1579_));
 sky130_fd_sc_hd__o21ai_2 _5591_ (.A1(_1578_),
    .A2(_1579_),
    .B1(\mul_la.reg_b0[13] ),
    .Y(_1580_));
 sky130_fd_sc_hd__or3_2 _5592_ (.A(\mul_la.reg_b0[13] ),
    .B(_1578_),
    .C(_1579_),
    .X(_1581_));
 sky130_fd_sc_hd__and2_2 _5593_ (.A(_1580_),
    .B(_1581_),
    .X(_1582_));
 sky130_fd_sc_hd__and3_1 _5594_ (.A(\mul_la.lob_4.L[2] ),
    .B(_1580_),
    .C(_1581_),
    .X(_1583_));
 sky130_fd_sc_hd__xor2_1 _5595_ (.A(\mul_la.reg_b0[13] ),
    .B(_1578_),
    .X(_1584_));
 sky130_fd_sc_hd__xnor2_4 _5596_ (.A(\mul_la.reg_b0[13] ),
    .B(_1578_),
    .Y(_1585_));
 sky130_fd_sc_hd__xor2_4 _5597_ (.A(\mul_la.reg_b0[12] ),
    .B(_1578_),
    .X(_1586_));
 sky130_fd_sc_hd__xnor2_4 _5598_ (.A(\mul_la.reg_b0[12] ),
    .B(_1578_),
    .Y(_1587_));
 sky130_fd_sc_hd__and3_1 _5599_ (.A(\mul_la.lob_4.L[3] ),
    .B(_1585_),
    .C(_1586_),
    .X(_1588_));
 sky130_fd_sc_hd__o21ba_1 _5600_ (.A1(_1583_),
    .A2(_1588_),
    .B1_N(_1577_),
    .X(_1589_));
 sky130_fd_sc_hd__o41a_4 _5601_ (.A1(_1565_),
    .A2(_1566_),
    .A3(_1567_),
    .A4(_1568_),
    .B1(net254),
    .X(_1590_));
 sky130_fd_sc_hd__and2_2 _5602_ (.A(net254),
    .B(\mul_la.reg_b0[10] ),
    .X(_1591_));
 sky130_fd_sc_hd__o21a_1 _5603_ (.A1(_1590_),
    .A2(_1591_),
    .B1(\mul_la.reg_b0[11] ),
    .X(_1592_));
 sky130_fd_sc_hd__o21ai_4 _5604_ (.A1(_1590_),
    .A2(_1591_),
    .B1(\mul_la.reg_b0[11] ),
    .Y(_1593_));
 sky130_fd_sc_hd__nor3_2 _5605_ (.A(\mul_la.reg_b0[11] ),
    .B(_1590_),
    .C(_1591_),
    .Y(_1594_));
 sky130_fd_sc_hd__or3_4 _5606_ (.A(\mul_la.reg_b0[11] ),
    .B(_1590_),
    .C(_1591_),
    .X(_1595_));
 sky130_fd_sc_hd__nor2_4 _5607_ (.A(_1592_),
    .B(_1594_),
    .Y(_1596_));
 sky130_fd_sc_hd__nand2_1 _5608_ (.A(_1593_),
    .B(_1595_),
    .Y(_1597_));
 sky130_fd_sc_hd__a21oi_4 _5609_ (.A1(_1593_),
    .A2(_1595_),
    .B1(_1586_),
    .Y(_1598_));
 sky130_fd_sc_hd__o211a_1 _5610_ (.A1(_3376_),
    .A2(_1573_),
    .B1(_1576_),
    .C1(_1585_),
    .X(_1599_));
 sky130_fd_sc_hd__xor2_4 _5611_ (.A(\mul_la.reg_b0[10] ),
    .B(_1590_),
    .X(_1600_));
 sky130_fd_sc_hd__xnor2_2 _5612_ (.A(\mul_la.reg_b0[10] ),
    .B(_1590_),
    .Y(_1601_));
 sky130_fd_sc_hd__o31a_2 _5613_ (.A1(_1565_),
    .A2(_1566_),
    .A3(_1567_),
    .B1(net254),
    .X(_1602_));
 sky130_fd_sc_hd__o41a_2 _5614_ (.A1(\mul_la.reg_b0[8] ),
    .A2(_1565_),
    .A3(_1566_),
    .A4(_1567_),
    .B1(net254),
    .X(_1603_));
 sky130_fd_sc_hd__xor2_4 _5615_ (.A(\mul_la.reg_b0[9] ),
    .B(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__xnor2_1 _5616_ (.A(\mul_la.reg_b0[9] ),
    .B(_1603_),
    .Y(_1605_));
 sky130_fd_sc_hd__and3_1 _5617_ (.A(\mul_la.lob_4.L[6] ),
    .B(_1601_),
    .C(_1604_),
    .X(_1606_));
 sky130_fd_sc_hd__and2_1 _5618_ (.A(\mul_la.lob_4.L[5] ),
    .B(_1600_),
    .X(_1607_));
 sky130_fd_sc_hd__xor2_4 _5619_ (.A(\mul_la.reg_b0[8] ),
    .B(_1602_),
    .X(_1608_));
 sky130_fd_sc_hd__and4_1 _5620_ (.A(\mul_la.lob_4.L[7] ),
    .B(_1601_),
    .C(_1605_),
    .D(_1608_),
    .X(_1609_));
 sky130_fd_sc_hd__o21a_2 _5621_ (.A1(_3376_),
    .A2(_1573_),
    .B1(_1575_),
    .X(_1610_));
 sky130_fd_sc_hd__o2111a_4 _5622_ (.A1(_3376_),
    .A2(_1573_),
    .B1(_1575_),
    .C1(_1585_),
    .D1(_1587_),
    .X(_1611_));
 sky130_fd_sc_hd__o211a_1 _5623_ (.A1(_1607_),
    .A2(_1609_),
    .B1(_1611_),
    .C1(_1597_),
    .X(_1612_));
 sky130_fd_sc_hd__a32o_1 _5624_ (.A1(_1598_),
    .A2(net235),
    .A3(_1606_),
    .B1(net236),
    .B2(\mul_la.lob_4.L[1] ),
    .X(_1613_));
 sky130_fd_sc_hd__nor3_1 _5625_ (.A(_1600_),
    .B(_1604_),
    .C(_1608_),
    .Y(_1614_));
 sky130_fd_sc_hd__o21a_1 _5626_ (.A1(_1565_),
    .A2(_1566_),
    .B1(net254),
    .X(_1615_));
 sky130_fd_sc_hd__o31a_4 _5627_ (.A1(\mul_la.reg_b0[6] ),
    .A2(_1565_),
    .A3(_1566_),
    .B1(net254),
    .X(_1616_));
 sky130_fd_sc_hd__xor2_4 _5628_ (.A(\mul_la.reg_b0[7] ),
    .B(_1616_),
    .X(_1617_));
 sky130_fd_sc_hd__xnor2_4 _5629_ (.A(\mul_la.reg_b0[7] ),
    .B(_1616_),
    .Y(_1618_));
 sky130_fd_sc_hd__nor4_2 _5630_ (.A(_1600_),
    .B(_1604_),
    .C(_1608_),
    .D(_1617_),
    .Y(_1619_));
 sky130_fd_sc_hd__and3_1 _5631_ (.A(_1598_),
    .B(net235),
    .C(_1619_),
    .X(_1620_));
 sky130_fd_sc_hd__xor2_4 _5632_ (.A(\mul_la.reg_b0[6] ),
    .B(_1615_),
    .X(_1621_));
 sky130_fd_sc_hd__o41a_2 _5633_ (.A1(\mul_la.reg_b0[1] ),
    .A2(\mul_la.lob_4.B[0] ),
    .A3(\mul_la.reg_b0[2] ),
    .A4(\mul_la.reg_b0[3] ),
    .B1(net254),
    .X(_1622_));
 sky130_fd_sc_hd__o211ai_2 _5634_ (.A1(\mul_la.reg_b0[4] ),
    .A2(_1565_),
    .B1(\mul_la.reg_b0[5] ),
    .C1(net254),
    .Y(_1623_));
 sky130_fd_sc_hd__a211o_1 _5635_ (.A1(net254),
    .A2(\mul_la.reg_b0[4] ),
    .B1(\mul_la.reg_b0[5] ),
    .C1(_1622_),
    .X(_1624_));
 sky130_fd_sc_hd__and2_2 _5636_ (.A(_1623_),
    .B(_1624_),
    .X(_1625_));
 sky130_fd_sc_hd__nand2_1 _5637_ (.A(_1623_),
    .B(_1624_),
    .Y(_1626_));
 sky130_fd_sc_hd__and3_1 _5638_ (.A(net264),
    .B(_1623_),
    .C(_1624_),
    .X(_1627_));
 sky130_fd_sc_hd__o31a_2 _5639_ (.A1(\mul_la.reg_b0[1] ),
    .A2(\mul_la.lob_4.B[0] ),
    .A3(\mul_la.reg_b0[2] ),
    .B1(net254),
    .X(_1628_));
 sky130_fd_sc_hd__xor2_4 _5640_ (.A(\mul_la.reg_b0[3] ),
    .B(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__xor2_4 _5641_ (.A(\mul_la.reg_b0[4] ),
    .B(_1622_),
    .X(_1630_));
 sky130_fd_sc_hd__nor2_2 _5642_ (.A(_1629_),
    .B(_1630_),
    .Y(_1631_));
 sky130_fd_sc_hd__o21ai_2 _5643_ (.A1(\mul_la.reg_b0[1] ),
    .A2(\mul_la.lob_4.B[0] ),
    .B1(net254),
    .Y(_1632_));
 sky130_fd_sc_hd__xnor2_4 _5644_ (.A(\mul_la.reg_b0[2] ),
    .B(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hd__nand2_2 _5645_ (.A(\mul_la.lob_4.B[0] ),
    .B(net254),
    .Y(_1634_));
 sky130_fd_sc_hd__xor2_2 _5646_ (.A(\mul_la.reg_b0[1] ),
    .B(_1634_),
    .X(_1635_));
 sky130_fd_sc_hd__xnor2_2 _5647_ (.A(\mul_la.reg_b0[1] ),
    .B(_1634_),
    .Y(_1636_));
 sky130_fd_sc_hd__nor2_1 _5648_ (.A(_1633_),
    .B(_1635_),
    .Y(_1637_));
 sky130_fd_sc_hd__and3_1 _5649_ (.A(_1626_),
    .B(_1631_),
    .C(_1637_),
    .X(_1638_));
 sky130_fd_sc_hd__a41o_1 _5650_ (.A1(net257),
    .A2(_1626_),
    .A3(_1631_),
    .A4(_1637_),
    .B1(_1627_),
    .X(_1639_));
 sky130_fd_sc_hd__nor2_1 _5651_ (.A(_1621_),
    .B(_1625_),
    .Y(_1640_));
 sky130_fd_sc_hd__nor2_1 _5652_ (.A(net236),
    .B(_1582_),
    .Y(_1641_));
 sky130_fd_sc_hd__and4_1 _5653_ (.A(\mul_la.lob_4.L[4] ),
    .B(\mul_la.lob_4.B[0] ),
    .C(_1587_),
    .D(_1596_),
    .X(_1642_));
 sky130_fd_sc_hd__and3_1 _5654_ (.A(\mul_la.lob_4.L[8] ),
    .B(\mul_la.lob_4.B[0] ),
    .C(_1617_),
    .X(_1643_));
 sky130_fd_sc_hd__and3_1 _5655_ (.A(_1598_),
    .B(_1614_),
    .C(_1643_),
    .X(_1644_));
 sky130_fd_sc_hd__o21a_1 _5656_ (.A1(_1642_),
    .A2(_1644_),
    .B1(_1641_),
    .X(_1645_));
 sky130_fd_sc_hd__a2111oi_4 _5657_ (.A1(_1593_),
    .A2(_1595_),
    .B1(_1600_),
    .C1(_1604_),
    .D1(_1608_),
    .Y(_1646_));
 sky130_fd_sc_hd__nor2_1 _5658_ (.A(_1617_),
    .B(_1621_),
    .Y(_1647_));
 sky130_fd_sc_hd__nor4_1 _5659_ (.A(_1584_),
    .B(_1586_),
    .C(_1617_),
    .D(_1621_),
    .Y(_1648_));
 sky130_fd_sc_hd__and2_1 _5660_ (.A(net234),
    .B(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__and4_1 _5661_ (.A(\mul_la.lob_4.B[0] ),
    .B(_1626_),
    .C(_1631_),
    .D(_1633_),
    .X(_1650_));
 sky130_fd_sc_hd__and4_1 _5662_ (.A(net259),
    .B(_1610_),
    .C(_1649_),
    .D(_1650_),
    .X(_1651_));
 sky130_fd_sc_hd__and2_1 _5663_ (.A(_1611_),
    .B(_1646_),
    .X(_1652_));
 sky130_fd_sc_hd__and4_1 _5664_ (.A(net265),
    .B(\mul_la.lob_4.B[0] ),
    .C(_1618_),
    .D(_1621_),
    .X(_1653_));
 sky130_fd_sc_hd__nor3_1 _5665_ (.A(_3372_),
    .B(_1633_),
    .C(_1636_),
    .Y(_1654_));
 sky130_fd_sc_hd__a22o_1 _5666_ (.A1(net263),
    .A2(_1630_),
    .B1(_1631_),
    .B2(_1654_),
    .X(_1655_));
 sky130_fd_sc_hd__a41o_1 _5667_ (.A1(\mul_la.lob_4.B[0] ),
    .A2(_1626_),
    .A3(_1647_),
    .A4(_1655_),
    .B1(_1653_),
    .X(_1656_));
 sky130_fd_sc_hd__o31a_1 _5668_ (.A1(_1589_),
    .A2(_1612_),
    .A3(_1613_),
    .B1(\mul_la.lob_4.B[0] ),
    .X(_1657_));
 sky130_fd_sc_hd__and3_1 _5669_ (.A(net261),
    .B(\mul_la.lob_4.B[0] ),
    .C(_1629_),
    .X(_1658_));
 sky130_fd_sc_hd__or4b_1 _5670_ (.A(_1621_),
    .B(_1625_),
    .C(_1630_),
    .D_N(_1658_),
    .X(_1659_));
 sky130_fd_sc_hd__and2b_1 _5671_ (.A_N(_1621_),
    .B(\mul_la.lob_4.B[0] ),
    .X(_1660_));
 sky130_fd_sc_hd__a21bo_1 _5672_ (.A1(_1639_),
    .A2(_1660_),
    .B1_N(_1659_),
    .X(_1661_));
 sky130_fd_sc_hd__a22o_1 _5673_ (.A1(_1652_),
    .A2(_1656_),
    .B1(_1661_),
    .B2(_1620_),
    .X(_1662_));
 sky130_fd_sc_hd__or4_2 _5674_ (.A(_1645_),
    .B(_1651_),
    .C(_1657_),
    .D(_1662_),
    .X(_1663_));
 sky130_fd_sc_hd__inv_2 _5675_ (.A(net188),
    .Y(_1664_));
 sky130_fd_sc_hd__or4_4 _5676_ (.A(\mul_la.reg_a0[2] ),
    .B(\mul_la.reg_a0[1] ),
    .C(\mul_la.lob_4.A[0] ),
    .D(\mul_la.reg_a0[3] ),
    .X(_1665_));
 sky130_fd_sc_hd__or2_4 _5677_ (.A(\mul_la.reg_a0[4] ),
    .B(\mul_la.reg_a0[5] ),
    .X(_1666_));
 sky130_fd_sc_hd__or2_2 _5678_ (.A(\mul_la.reg_a0[6] ),
    .B(\mul_la.reg_a0[7] ),
    .X(_1667_));
 sky130_fd_sc_hd__o31a_1 _5679_ (.A1(_1665_),
    .A2(_1666_),
    .A3(_1667_),
    .B1(net253),
    .X(_1668_));
 sky130_fd_sc_hd__o41a_2 _5680_ (.A1(\mul_la.reg_a0[8] ),
    .A2(_1665_),
    .A3(_1666_),
    .A4(_1667_),
    .B1(net253),
    .X(_1669_));
 sky130_fd_sc_hd__xor2_4 _5681_ (.A(\mul_la.reg_a0[9] ),
    .B(_1669_),
    .X(_1670_));
 sky130_fd_sc_hd__o31a_1 _5682_ (.A1(_1665_),
    .A2(_1666_),
    .A3(_1667_),
    .B1(\mul_la.reg_a0[8] ),
    .X(_1671_));
 sky130_fd_sc_hd__o2bb2a_4 _5683_ (.A1_N(net253),
    .A2_N(_1671_),
    .B1(_1668_),
    .B2(\mul_la.reg_a0[8] ),
    .X(_1672_));
 sky130_fd_sc_hd__or2_1 _5684_ (.A(\mul_la.reg_a0[8] ),
    .B(\mul_la.reg_a0[9] ),
    .X(_1673_));
 sky130_fd_sc_hd__o41a_4 _5685_ (.A1(_1665_),
    .A2(_1666_),
    .A3(_1667_),
    .A4(_1673_),
    .B1(net253),
    .X(_1674_));
 sky130_fd_sc_hd__xnor2_4 _5686_ (.A(\mul_la.reg_a0[10] ),
    .B(_1674_),
    .Y(_1675_));
 sky130_fd_sc_hd__xor2_4 _5687_ (.A(\mul_la.reg_a0[10] ),
    .B(_1674_),
    .X(_1676_));
 sky130_fd_sc_hd__and2_1 _5688_ (.A(net253),
    .B(\mul_la.reg_a0[10] ),
    .X(_1677_));
 sky130_fd_sc_hd__o21ai_4 _5689_ (.A1(_1674_),
    .A2(_1677_),
    .B1(\mul_la.reg_a0[11] ),
    .Y(_1678_));
 sky130_fd_sc_hd__or3_4 _5690_ (.A(\mul_la.reg_a0[11] ),
    .B(_1674_),
    .C(_1677_),
    .X(_1679_));
 sky130_fd_sc_hd__and2_4 _5691_ (.A(_1678_),
    .B(_1679_),
    .X(_1680_));
 sky130_fd_sc_hd__a21oi_4 _5692_ (.A1(_1678_),
    .A2(_1679_),
    .B1(_1676_),
    .Y(_1681_));
 sky130_fd_sc_hd__or4_1 _5693_ (.A(\mul_la.reg_a0[8] ),
    .B(\mul_la.reg_a0[9] ),
    .C(\mul_la.reg_a0[10] ),
    .D(\mul_la.reg_a0[11] ),
    .X(_1682_));
 sky130_fd_sc_hd__or4_2 _5694_ (.A(_1665_),
    .B(_1666_),
    .C(_1667_),
    .D(_1682_),
    .X(_1683_));
 sky130_fd_sc_hd__o21a_2 _5695_ (.A1(\mul_la.reg_a0[12] ),
    .A2(_1683_),
    .B1(net253),
    .X(_1684_));
 sky130_fd_sc_hd__xor2_4 _5696_ (.A(\mul_la.reg_a0[13] ),
    .B(_1684_),
    .X(_1685_));
 sky130_fd_sc_hd__xnor2_4 _5697_ (.A(\mul_la.reg_a0[13] ),
    .B(_1684_),
    .Y(_1686_));
 sky130_fd_sc_hd__o41a_2 _5698_ (.A1(_1665_),
    .A2(_1666_),
    .A3(_1667_),
    .A4(_1682_),
    .B1(net253),
    .X(_1687_));
 sky130_fd_sc_hd__xor2_4 _5699_ (.A(\mul_la.reg_a0[12] ),
    .B(_1687_),
    .X(_1688_));
 sky130_fd_sc_hd__nor2_1 _5700_ (.A(_1685_),
    .B(_1688_),
    .Y(_1689_));
 sky130_fd_sc_hd__nor2_1 _5701_ (.A(\mul_la.reg_a0[12] ),
    .B(\mul_la.reg_a0[13] ),
    .Y(_1690_));
 sky130_fd_sc_hd__o31a_2 _5702_ (.A1(\mul_la.reg_a0[12] ),
    .A2(\mul_la.reg_a0[13] ),
    .A3(_1683_),
    .B1(net253),
    .X(_1691_));
 sky130_fd_sc_hd__xnor2_2 _5703_ (.A(\mul_la.reg_a0[14] ),
    .B(_1691_),
    .Y(_1692_));
 sky130_fd_sc_hd__xor2_4 _5704_ (.A(\mul_la.reg_a0[14] ),
    .B(_1691_),
    .X(_1693_));
 sky130_fd_sc_hd__and4bb_4 _5705_ (.A_N(\mul_la.reg_a0[14] ),
    .B_N(_1683_),
    .C(_1690_),
    .D(net253),
    .X(_1694_));
 sky130_fd_sc_hd__nor2_2 _5706_ (.A(net232),
    .B(_1694_),
    .Y(_1695_));
 sky130_fd_sc_hd__nor4_4 _5707_ (.A(_1685_),
    .B(_1688_),
    .C(net232),
    .D(_1694_),
    .Y(_1696_));
 sky130_fd_sc_hd__o21ai_4 _5708_ (.A1(_1665_),
    .A2(_1666_),
    .B1(net253),
    .Y(_1697_));
 sky130_fd_sc_hd__o31a_2 _5709_ (.A1(\mul_la.reg_a0[6] ),
    .A2(_1665_),
    .A3(_1666_),
    .B1(net253),
    .X(_1698_));
 sky130_fd_sc_hd__xor2_4 _5710_ (.A(\mul_la.reg_a0[7] ),
    .B(_1698_),
    .X(_1699_));
 sky130_fd_sc_hd__xnor2_4 _5711_ (.A(\mul_la.reg_a0[6] ),
    .B(_1697_),
    .Y(_1700_));
 sky130_fd_sc_hd__and3b_1 _5712_ (.A_N(_1699_),
    .B(_1696_),
    .C(_1681_),
    .X(_1701_));
 sky130_fd_sc_hd__nand2_2 _5713_ (.A(_1686_),
    .B(net233),
    .Y(_1702_));
 sky130_fd_sc_hd__a21oi_4 _5714_ (.A1(_1678_),
    .A2(_1679_),
    .B1(_1688_),
    .Y(_1703_));
 sky130_fd_sc_hd__and3_2 _5715_ (.A(_1686_),
    .B(net233),
    .C(_1703_),
    .X(_1704_));
 sky130_fd_sc_hd__and4_1 _5716_ (.A(\mul_la.lob_4.L[8] ),
    .B(_1675_),
    .C(_1699_),
    .D(_1704_),
    .X(_1705_));
 sky130_fd_sc_hd__a31o_1 _5717_ (.A1(net265),
    .A2(_1700_),
    .A3(_1701_),
    .B1(_1705_),
    .X(_1706_));
 sky130_fd_sc_hd__o41a_2 _5718_ (.A1(\mul_la.reg_a0[2] ),
    .A2(\mul_la.reg_a0[1] ),
    .A3(\mul_la.lob_4.A[0] ),
    .A4(\mul_la.reg_a0[3] ),
    .B1(net253),
    .X(_1707_));
 sky130_fd_sc_hd__a21oi_2 _5719_ (.A1(net253),
    .A2(\mul_la.reg_a0[4] ),
    .B1(_1707_),
    .Y(_1708_));
 sky130_fd_sc_hd__xnor2_4 _5720_ (.A(\mul_la.reg_a0[5] ),
    .B(_1708_),
    .Y(_1709_));
 sky130_fd_sc_hd__or2_1 _5721_ (.A(_1700_),
    .B(_1709_),
    .X(_1710_));
 sky130_fd_sc_hd__nor2_1 _5722_ (.A(_1670_),
    .B(_1676_),
    .Y(_1711_));
 sky130_fd_sc_hd__nor2_1 _5723_ (.A(_1672_),
    .B(_1699_),
    .Y(_1712_));
 sky130_fd_sc_hd__nor4_1 _5724_ (.A(_1670_),
    .B(_1672_),
    .C(_1676_),
    .D(_1699_),
    .Y(_1713_));
 sky130_fd_sc_hd__or4_1 _5725_ (.A(_1670_),
    .B(_1672_),
    .C(_1676_),
    .D(_1699_),
    .X(_1714_));
 sky130_fd_sc_hd__and4_2 _5726_ (.A(_1686_),
    .B(net233),
    .C(_1703_),
    .D(_1713_),
    .X(_1715_));
 sky130_fd_sc_hd__o21ai_2 _5727_ (.A1(\mul_la.reg_a0[1] ),
    .A2(\mul_la.lob_4.A[0] ),
    .B1(net253),
    .Y(_1716_));
 sky130_fd_sc_hd__o31a_2 _5728_ (.A1(\mul_la.reg_a0[2] ),
    .A2(\mul_la.reg_a0[1] ),
    .A3(\mul_la.lob_4.A[0] ),
    .B1(net253),
    .X(_1717_));
 sky130_fd_sc_hd__xor2_1 _5729_ (.A(\mul_la.reg_a0[3] ),
    .B(_1717_),
    .X(_1718_));
 sky130_fd_sc_hd__xnor2_4 _5730_ (.A(\mul_la.reg_a0[3] ),
    .B(_1717_),
    .Y(_1719_));
 sky130_fd_sc_hd__xor2_4 _5731_ (.A(\mul_la.reg_a0[4] ),
    .B(_1707_),
    .X(_1720_));
 sky130_fd_sc_hd__nor2_1 _5732_ (.A(_1718_),
    .B(_1720_),
    .Y(_1721_));
 sky130_fd_sc_hd__xor2_1 _5733_ (.A(\mul_la.reg_a0[2] ),
    .B(_1716_),
    .X(_1722_));
 sky130_fd_sc_hd__xnor2_1 _5734_ (.A(\mul_la.reg_a0[2] ),
    .B(_1716_),
    .Y(_1723_));
 sky130_fd_sc_hd__nand2_2 _5735_ (.A(\mul_la.lob_4.A[0] ),
    .B(net253),
    .Y(_1724_));
 sky130_fd_sc_hd__xor2_4 _5736_ (.A(\mul_la.reg_a0[1] ),
    .B(_1724_),
    .X(_1725_));
 sky130_fd_sc_hd__nor2_1 _5737_ (.A(_1670_),
    .B(_1672_),
    .Y(_1726_));
 sky130_fd_sc_hd__a2111oi_2 _5738_ (.A1(_1678_),
    .A2(_1679_),
    .B1(_1670_),
    .C1(_1672_),
    .D1(_1676_),
    .Y(_1727_));
 sky130_fd_sc_hd__nor3_1 _5739_ (.A(_1718_),
    .B(_1720_),
    .C(_1722_),
    .Y(_1728_));
 sky130_fd_sc_hd__a22o_1 _5740_ (.A1(net263),
    .A2(_1720_),
    .B1(_1728_),
    .B2(net259),
    .X(_1729_));
 sky130_fd_sc_hd__nor2_1 _5741_ (.A(_1699_),
    .B(_1700_),
    .Y(_1730_));
 sky130_fd_sc_hd__and4bb_2 _5742_ (.A_N(_1685_),
    .B_N(_1688_),
    .C(_1727_),
    .D(_1730_),
    .X(_1731_));
 sky130_fd_sc_hd__or3_4 _5743_ (.A(_3372_),
    .B(net232),
    .C(_1694_),
    .X(_1732_));
 sky130_fd_sc_hd__nor4b_4 _5744_ (.A(_1709_),
    .B(_1732_),
    .C(_1720_),
    .D_N(_1731_),
    .Y(_1733_));
 sky130_fd_sc_hd__and3_1 _5745_ (.A(_1719_),
    .B(_1722_),
    .C(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__and4_1 _5746_ (.A(\mul_la.lob_4.L[6] ),
    .B(_1670_),
    .C(_1675_),
    .D(_1704_),
    .X(_1735_));
 sky130_fd_sc_hd__a21oi_1 _5747_ (.A1(_1678_),
    .A2(_1679_),
    .B1(_1675_),
    .Y(_1736_));
 sky130_fd_sc_hd__a221o_1 _5748_ (.A1(\mul_la.lob_4.L[4] ),
    .A2(_1680_),
    .B1(_1736_),
    .B2(\mul_la.lob_4.L[5] ),
    .C1(_1688_),
    .X(_1737_));
 sky130_fd_sc_hd__a211oi_1 _5749_ (.A1(_3375_),
    .A2(_1688_),
    .B1(net232),
    .C1(_1685_),
    .Y(_1738_));
 sky130_fd_sc_hd__and2_1 _5750_ (.A(\mul_la.lob_4.L[1] ),
    .B(net232),
    .X(_1739_));
 sky130_fd_sc_hd__nor2_2 _5751_ (.A(_1686_),
    .B(net232),
    .Y(_1740_));
 sky130_fd_sc_hd__nand2_2 _5752_ (.A(_1685_),
    .B(net233),
    .Y(_1741_));
 sky130_fd_sc_hd__and3_1 _5753_ (.A(\mul_la.lob_4.L[2] ),
    .B(_1685_),
    .C(_1692_),
    .X(_1742_));
 sky130_fd_sc_hd__a211o_1 _5754_ (.A1(_1737_),
    .A2(_1738_),
    .B1(_1739_),
    .C1(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__nor3_1 _5755_ (.A(_1709_),
    .B(_1719_),
    .C(_1720_),
    .Y(_1744_));
 sky130_fd_sc_hd__a22o_1 _5756_ (.A1(net264),
    .A2(_1709_),
    .B1(_1744_),
    .B2(net261),
    .X(_1745_));
 sky130_fd_sc_hd__and3b_1 _5757_ (.A_N(_1700_),
    .B(_1715_),
    .C(_1745_),
    .X(_1746_));
 sky130_fd_sc_hd__and3b_1 _5758_ (.A_N(_1670_),
    .B(_1672_),
    .C(\mul_la.lob_4.L[7] ),
    .X(_1747_));
 sky130_fd_sc_hd__and3_1 _5759_ (.A(_1681_),
    .B(net226),
    .C(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__or4_1 _5760_ (.A(_1735_),
    .B(_1743_),
    .C(_1746_),
    .D(_1748_),
    .X(_1749_));
 sky130_fd_sc_hd__a221o_1 _5761_ (.A1(_1706_),
    .A2(_1726_),
    .B1(_1734_),
    .B2(_1725_),
    .C1(_1749_),
    .X(_1750_));
 sky130_fd_sc_hd__and4b_1 _5762_ (.A_N(_1725_),
    .B(_1722_),
    .C(net257),
    .D(\mul_la.lob_4.A[0] ),
    .X(_1751_));
 sky130_fd_sc_hd__and3b_1 _5763_ (.A_N(_1699_),
    .B(_1729_),
    .C(\mul_la.lob_4.A[0] ),
    .X(_1752_));
 sky130_fd_sc_hd__and3_1 _5764_ (.A(_1696_),
    .B(_1727_),
    .C(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__a31oi_1 _5765_ (.A1(_1715_),
    .A2(_1721_),
    .A3(_1751_),
    .B1(_1753_),
    .Y(_1754_));
 sky130_fd_sc_hd__o2bb2a_4 _5766_ (.A1_N(net709),
    .A2_N(_1750_),
    .B1(_1754_),
    .B2(_1710_),
    .X(_1755_));
 sky130_fd_sc_hd__inv_2 _5767_ (.A(_1755_),
    .Y(_1756_));
 sky130_fd_sc_hd__nor2_2 _5768_ (.A(_1664_),
    .B(_1755_),
    .Y(\mul_la.P_[0] ));
 sky130_fd_sc_hd__and3_4 _5769_ (.A(_1696_),
    .B(_1699_),
    .C(_1727_),
    .X(_1757_));
 sky130_fd_sc_hd__nor2_1 _5770_ (.A(_1710_),
    .B(_1714_),
    .Y(_1758_));
 sky130_fd_sc_hd__a22o_1 _5771_ (.A1(net261),
    .A2(_1720_),
    .B1(_1728_),
    .B2(net257),
    .X(_1759_));
 sky130_fd_sc_hd__and3b_1 _5772_ (.A_N(_1710_),
    .B(_1713_),
    .C(_1759_),
    .X(_1760_));
 sky130_fd_sc_hd__and3b_1 _5773_ (.A_N(_1670_),
    .B(_1672_),
    .C(_1675_),
    .X(_1761_));
 sky130_fd_sc_hd__a22o_1 _5774_ (.A1(\mul_la.lob_4.L[6] ),
    .A2(_1676_),
    .B1(_1761_),
    .B2(\mul_la.lob_4.L[8] ),
    .X(_1762_));
 sky130_fd_sc_hd__o21ai_1 _5775_ (.A1(_1760_),
    .A2(_1762_),
    .B1(_1703_),
    .Y(_1763_));
 sky130_fd_sc_hd__a21boi_1 _5776_ (.A1(\mul_la.lob_4.L[4] ),
    .A2(_1688_),
    .B1_N(_1763_),
    .Y(_1764_));
 sky130_fd_sc_hd__a32o_1 _5777_ (.A1(net264),
    .A2(_1700_),
    .A3(_1715_),
    .B1(_1757_),
    .B2(net265),
    .X(_1765_));
 sky130_fd_sc_hd__o21ba_2 _5778_ (.A1(_1702_),
    .A2(_1764_),
    .B1_N(_1765_),
    .X(_1766_));
 sky130_fd_sc_hd__a22o_1 _5779_ (.A1(\mul_la.lob_4.L[2] ),
    .A2(_1693_),
    .B1(_1740_),
    .B2(\mul_la.lob_4.L[3] ),
    .X(_1767_));
 sky130_fd_sc_hd__and2_1 _5780_ (.A(_1680_),
    .B(net226),
    .X(_1768_));
 sky130_fd_sc_hd__and3b_1 _5781_ (.A_N(_1694_),
    .B(_1709_),
    .C(_1692_),
    .X(_1769_));
 sky130_fd_sc_hd__and3_1 _5782_ (.A(net263),
    .B(_1731_),
    .C(_1769_),
    .X(_1770_));
 sky130_fd_sc_hd__and4_1 _5783_ (.A(net259),
    .B(_1695_),
    .C(_1731_),
    .D(_1744_),
    .X(_1771_));
 sky130_fd_sc_hd__a2111o_1 _5784_ (.A1(\mul_la.lob_4.L[5] ),
    .A2(_1768_),
    .B1(_1770_),
    .C1(_1771_),
    .D1(_1767_),
    .X(_1772_));
 sky130_fd_sc_hd__and3_4 _5785_ (.A(_1670_),
    .B(_1681_),
    .C(net226),
    .X(_1773_));
 sky130_fd_sc_hd__a211oi_4 _5786_ (.A1(\mul_la.lob_4.L[7] ),
    .A2(_1773_),
    .B1(_1772_),
    .C1(_1734_),
    .Y(_1774_));
 sky130_fd_sc_hd__a21oi_2 _5787_ (.A1(_1766_),
    .A2(_1774_),
    .B1(_1725_),
    .Y(_1775_));
 sky130_fd_sc_hd__a21o_2 _5788_ (.A1(_1766_),
    .A2(_1774_),
    .B1(_1725_),
    .X(_1776_));
 sky130_fd_sc_hd__and3_1 _5789_ (.A(_1611_),
    .B(_1617_),
    .C(net234),
    .X(_1777_));
 sky130_fd_sc_hd__and4_1 _5790_ (.A(net265),
    .B(_1611_),
    .C(_1617_),
    .D(_1646_),
    .X(_1778_));
 sky130_fd_sc_hd__and3_1 _5791_ (.A(_1598_),
    .B(net235),
    .C(_1600_),
    .X(_1779_));
 sky130_fd_sc_hd__and4_1 _5792_ (.A(\mul_la.lob_4.L[6] ),
    .B(_1598_),
    .C(_1599_),
    .D(_1600_),
    .X(_1780_));
 sky130_fd_sc_hd__o2111a_2 _5793_ (.A1(_1592_),
    .A2(_1594_),
    .B1(_1601_),
    .C1(_1587_),
    .D1(_1585_),
    .X(_1781_));
 sky130_fd_sc_hd__o211a_2 _5794_ (.A1(_3376_),
    .A2(_1573_),
    .B1(_1575_),
    .C1(_1604_),
    .X(_1782_));
 sky130_fd_sc_hd__and3_1 _5795_ (.A(\mul_la.lob_4.L[7] ),
    .B(_1781_),
    .C(_1782_),
    .X(_1783_));
 sky130_fd_sc_hd__o2111a_4 _5796_ (.A1(_3376_),
    .A2(_1573_),
    .B1(_1575_),
    .C1(_1580_),
    .D1(_1581_),
    .X(_1784_));
 sky130_fd_sc_hd__a22o_1 _5797_ (.A1(\mul_la.lob_4.L[2] ),
    .A2(net236),
    .B1(_1784_),
    .B2(\mul_la.lob_4.L[3] ),
    .X(_1785_));
 sky130_fd_sc_hd__nor4_1 _5798_ (.A(_1778_),
    .B(_1780_),
    .C(_1783_),
    .D(_1785_),
    .Y(_1786_));
 sky130_fd_sc_hd__and4_2 _5799_ (.A(_1598_),
    .B(net235),
    .C(_1619_),
    .D(_1621_),
    .X(_1787_));
 sky130_fd_sc_hd__nand2_1 _5800_ (.A(net264),
    .B(_1787_),
    .Y(_1788_));
 sky130_fd_sc_hd__o2111a_2 _5801_ (.A1(_1592_),
    .A2(_1594_),
    .B1(_1601_),
    .C1(_1605_),
    .D1(_1587_),
    .X(_1789_));
 sky130_fd_sc_hd__a32o_1 _5802_ (.A1(net258),
    .A2(_1631_),
    .A3(_1633_),
    .B1(net261),
    .B2(_1630_),
    .X(_1790_));
 sky130_fd_sc_hd__and4_1 _5803_ (.A(_1598_),
    .B(_1619_),
    .C(_1640_),
    .D(_1790_),
    .X(_1791_));
 sky130_fd_sc_hd__a32o_1 _5804_ (.A1(\mul_la.lob_4.L[8] ),
    .A2(_1608_),
    .A3(_1789_),
    .B1(\mul_la.lob_4.L[4] ),
    .B2(_1586_),
    .X(_1792_));
 sky130_fd_sc_hd__o21ai_1 _5805_ (.A1(_1791_),
    .A2(_1792_),
    .B1(net235),
    .Y(_1793_));
 sky130_fd_sc_hd__a31o_4 _5806_ (.A1(_1786_),
    .A2(_1788_),
    .A3(_1793_),
    .B1(_1635_),
    .X(_1794_));
 sky130_fd_sc_hd__and3_1 _5807_ (.A(net256),
    .B(_1610_),
    .C(_1638_),
    .X(_1795_));
 sky130_fd_sc_hd__o211a_1 _5808_ (.A1(_3376_),
    .A2(_1573_),
    .B1(_1575_),
    .C1(_1625_),
    .X(_1796_));
 sky130_fd_sc_hd__a31o_1 _5809_ (.A1(\mul_la.lob_4.L[11] ),
    .A2(_1636_),
    .A3(_1796_),
    .B1(_1795_),
    .X(_1797_));
 sky130_fd_sc_hd__and2_1 _5810_ (.A(_1596_),
    .B(_1611_),
    .X(_1798_));
 sky130_fd_sc_hd__nor4_1 _5811_ (.A(_1617_),
    .B(_1621_),
    .C(_1625_),
    .D(_1630_),
    .Y(_1799_));
 sky130_fd_sc_hd__and4_1 _5812_ (.A(net259),
    .B(_1629_),
    .C(_1636_),
    .D(_1799_),
    .X(_1800_));
 sky130_fd_sc_hd__a32o_1 _5813_ (.A1(\mul_la.lob_4.L[5] ),
    .A2(_1636_),
    .A3(_1798_),
    .B1(_1800_),
    .B2(_1652_),
    .X(_1801_));
 sky130_fd_sc_hd__a21oi_4 _5814_ (.A1(_1649_),
    .A2(_1797_),
    .B1(_1801_),
    .Y(_1802_));
 sky130_fd_sc_hd__and2_1 _5815_ (.A(_1794_),
    .B(_1802_),
    .X(_1803_));
 sky130_fd_sc_hd__nand2_4 _5816_ (.A(_1794_),
    .B(_1802_),
    .Y(_1804_));
 sky130_fd_sc_hd__a22o_1 _5817_ (.A1(net188),
    .A2(net167),
    .B1(_1804_),
    .B2(_1756_),
    .X(_1805_));
 sky130_fd_sc_hd__inv_2 _5818_ (.A(_1805_),
    .Y(_1806_));
 sky130_fd_sc_hd__and4_1 _5819_ (.A(net188),
    .B(_1756_),
    .C(net167),
    .D(_1804_),
    .X(_1807_));
 sky130_fd_sc_hd__xor2_1 _5820_ (.A(\mul_la.reg_a0[15] ),
    .B(net699),
    .X(_1808_));
 sky130_fd_sc_hd__xnor2_4 _5821_ (.A(net704),
    .B(net699),
    .Y(_1809_));
 sky130_fd_sc_hd__o211ai_1 _5822_ (.A1(_1806_),
    .A2(_1807_),
    .B1(net251),
    .C1(\mul_la.P_[0] ),
    .Y(_1810_));
 sky130_fd_sc_hd__a211o_1 _5823_ (.A1(\mul_la.P_[0] ),
    .A2(net251),
    .B1(_1807_),
    .C1(_1806_),
    .X(_1811_));
 sky130_fd_sc_hd__nand2_1 _5824_ (.A(_1810_),
    .B(_1811_),
    .Y(\mul_la.reg_p[1] ));
 sky130_fd_sc_hd__and3_1 _5825_ (.A(net235),
    .B(_1608_),
    .C(_1789_),
    .X(_1812_));
 sky130_fd_sc_hd__and2_1 _5826_ (.A(net264),
    .B(_1777_),
    .X(_1813_));
 sky130_fd_sc_hd__a32o_1 _5827_ (.A1(net263),
    .A2(_1619_),
    .A3(_1621_),
    .B1(\mul_la.lob_4.L[7] ),
    .B2(_1600_),
    .X(_1814_));
 sky130_fd_sc_hd__and3_1 _5828_ (.A(\mul_la.lob_4.L[6] ),
    .B(_1593_),
    .C(_1595_),
    .X(_1815_));
 sky130_fd_sc_hd__a41o_1 _5829_ (.A1(\mul_la.lob_4.L[8] ),
    .A2(_1597_),
    .A3(_1601_),
    .A4(_1604_),
    .B1(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__a32o_1 _5830_ (.A1(_1585_),
    .A2(_1587_),
    .A3(_1816_),
    .B1(_1582_),
    .B2(\mul_la.lob_4.L[4] ),
    .X(_1817_));
 sky130_fd_sc_hd__o2111a_4 _5831_ (.A1(_3376_),
    .A2(_1573_),
    .B1(_1576_),
    .C1(_1585_),
    .D1(_1586_),
    .X(_1818_));
 sky130_fd_sc_hd__a22o_1 _5832_ (.A1(\mul_la.lob_4.L[3] ),
    .A2(_1577_),
    .B1(_1818_),
    .B2(\mul_la.lob_4.L[5] ),
    .X(_1819_));
 sky130_fd_sc_hd__and3_1 _5833_ (.A(net258),
    .B(_1611_),
    .C(_1629_),
    .X(_1820_));
 sky130_fd_sc_hd__and3_1 _5834_ (.A(net234),
    .B(net231),
    .C(_1820_),
    .X(_1821_));
 sky130_fd_sc_hd__and4_1 _5835_ (.A(_1598_),
    .B(net235),
    .C(_1619_),
    .D(_1640_),
    .X(_1822_));
 sky130_fd_sc_hd__and3_1 _5836_ (.A(net255),
    .B(_1631_),
    .C(_1822_),
    .X(_1823_));
 sky130_fd_sc_hd__a32o_1 _5837_ (.A1(_1598_),
    .A2(net235),
    .A3(_1814_),
    .B1(_1812_),
    .B2(net265),
    .X(_1824_));
 sky130_fd_sc_hd__a311o_1 _5838_ (.A1(net261),
    .A2(_1649_),
    .A3(_1796_),
    .B1(_1821_),
    .C1(_1824_),
    .X(_1825_));
 sky130_fd_sc_hd__and3_1 _5839_ (.A(net259),
    .B(_1630_),
    .C(_1822_),
    .X(_1826_));
 sky130_fd_sc_hd__a211o_1 _5840_ (.A1(_1610_),
    .A2(_1817_),
    .B1(_1823_),
    .C1(_1826_),
    .X(_1827_));
 sky130_fd_sc_hd__o41a_2 _5841_ (.A1(_1813_),
    .A2(_1819_),
    .A3(_1825_),
    .A4(_1827_),
    .B1(_1633_),
    .X(_1828_));
 sky130_fd_sc_hd__o41ai_4 _5842_ (.A1(_1813_),
    .A2(_1819_),
    .A3(_1825_),
    .A4(_1827_),
    .B1(_1633_),
    .Y(_1829_));
 sky130_fd_sc_hd__nor2_1 _5843_ (.A(_1755_),
    .B(_1829_),
    .Y(_1830_));
 sky130_fd_sc_hd__nand2_1 _5844_ (.A(net167),
    .B(_1804_),
    .Y(_1831_));
 sky130_fd_sc_hd__or4b_1 _5845_ (.A(_3373_),
    .B(_1710_),
    .C(_1714_),
    .D_N(_1720_),
    .X(_1832_));
 sky130_fd_sc_hd__nand2_1 _5846_ (.A(\mul_la.lob_4.L[7] ),
    .B(_1676_),
    .Y(_1833_));
 sky130_fd_sc_hd__a32o_1 _5847_ (.A1(net263),
    .A2(_1700_),
    .A3(_1712_),
    .B1(net265),
    .B2(_1672_),
    .X(_1834_));
 sky130_fd_sc_hd__and3_2 _5848_ (.A(_1686_),
    .B(_1688_),
    .C(net233),
    .X(_1835_));
 sky130_fd_sc_hd__a22o_1 _5849_ (.A1(\mul_la.lob_4.L[3] ),
    .A2(net232),
    .B1(_1835_),
    .B2(\mul_la.lob_4.L[5] ),
    .X(_1836_));
 sky130_fd_sc_hd__and4_1 _5850_ (.A(net257),
    .B(_1695_),
    .C(_1731_),
    .D(_1744_),
    .X(_1837_));
 sky130_fd_sc_hd__a32o_1 _5851_ (.A1(\mul_la.lob_4.L[6] ),
    .A2(_1680_),
    .A3(_1689_),
    .B1(_1685_),
    .B2(\mul_la.lob_4.L[4] ),
    .X(_1838_));
 sky130_fd_sc_hd__and4_1 _5852_ (.A(net256),
    .B(_1686_),
    .C(net233),
    .D(_1703_),
    .X(_1839_));
 sky130_fd_sc_hd__and3_1 _5853_ (.A(_1721_),
    .B(_1758_),
    .C(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__a21boi_1 _5854_ (.A1(_1832_),
    .A2(_1833_),
    .B1_N(_1704_),
    .Y(_1841_));
 sky130_fd_sc_hd__and3_1 _5855_ (.A(_1704_),
    .B(_1711_),
    .C(_1834_),
    .X(_1842_));
 sky130_fd_sc_hd__and3_1 _5856_ (.A(net261),
    .B(_1731_),
    .C(_1769_),
    .X(_1843_));
 sky130_fd_sc_hd__or4_1 _5857_ (.A(_1837_),
    .B(_1841_),
    .C(_1842_),
    .D(_1843_),
    .X(_1844_));
 sky130_fd_sc_hd__a211o_1 _5858_ (.A1(_1695_),
    .A2(_1838_),
    .B1(_1840_),
    .C1(_1836_),
    .X(_1845_));
 sky130_fd_sc_hd__a22o_1 _5859_ (.A1(net264),
    .A2(_1757_),
    .B1(_1773_),
    .B2(\mul_la.lob_4.L[8] ),
    .X(_1846_));
 sky130_fd_sc_hd__o31ai_1 _5860_ (.A1(_1844_),
    .A2(_1845_),
    .A3(_1846_),
    .B1(_1723_),
    .Y(_1847_));
 sky130_fd_sc_hd__nor2_1 _5861_ (.A(_1664_),
    .B(net170),
    .Y(_1848_));
 sky130_fd_sc_hd__xnor2_1 _5862_ (.A(_1831_),
    .B(_1848_),
    .Y(_1849_));
 sky130_fd_sc_hd__xor2_1 _5863_ (.A(_1830_),
    .B(_1849_),
    .X(_1850_));
 sky130_fd_sc_hd__nand2_1 _5864_ (.A(_1807_),
    .B(_1850_),
    .Y(_1851_));
 sky130_fd_sc_hd__or2_1 _5865_ (.A(_1807_),
    .B(_1850_),
    .X(_1852_));
 sky130_fd_sc_hd__nand2_1 _5866_ (.A(_1851_),
    .B(_1852_),
    .Y(_1853_));
 sky130_fd_sc_hd__o21ba_1 _5867_ (.A1(\mul_la.P_[0] ),
    .A2(_1805_),
    .B1_N(_1853_),
    .X(_1854_));
 sky130_fd_sc_hd__or3_1 _5868_ (.A(\mul_la.P_[0] ),
    .B(_1805_),
    .C(_1850_),
    .X(_1855_));
 sky130_fd_sc_hd__nand2_1 _5869_ (.A(net251),
    .B(_1855_),
    .Y(_1856_));
 sky130_fd_sc_hd__o22ai_1 _5870_ (.A1(net251),
    .A2(_1853_),
    .B1(_1854_),
    .B2(_1856_),
    .Y(\mul_la.reg_p[2] ));
 sky130_fd_sc_hd__a32o_1 _5871_ (.A1(net255),
    .A2(net234),
    .A3(net231),
    .B1(\mul_la.lob_4.L[7] ),
    .B2(_1596_),
    .X(_1857_));
 sky130_fd_sc_hd__and2_1 _5872_ (.A(_1611_),
    .B(_1857_),
    .X(_1858_));
 sky130_fd_sc_hd__and2_1 _5873_ (.A(\mul_la.lob_4.L[6] ),
    .B(_1818_),
    .X(_1859_));
 sky130_fd_sc_hd__and3_1 _5874_ (.A(net265),
    .B(_1781_),
    .C(_1782_),
    .X(_1860_));
 sky130_fd_sc_hd__and2_1 _5875_ (.A(\mul_la.lob_4.L[5] ),
    .B(_1784_),
    .X(_1861_));
 sky130_fd_sc_hd__a22o_1 _5876_ (.A1(\mul_la.lob_4.L[4] ),
    .A2(_1577_),
    .B1(_1784_),
    .B2(\mul_la.lob_4.L[5] ),
    .X(_1862_));
 sky130_fd_sc_hd__a2111o_1 _5877_ (.A1(net261),
    .A2(_1787_),
    .B1(_1859_),
    .C1(_1860_),
    .D1(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__and3_1 _5878_ (.A(net258),
    .B(_1630_),
    .C(_1822_),
    .X(_1864_));
 sky130_fd_sc_hd__and4_1 _5879_ (.A(net263),
    .B(_1611_),
    .C(_1617_),
    .D(net234),
    .X(_1865_));
 sky130_fd_sc_hd__and4_1 _5880_ (.A(\mul_la.lob_4.L[8] ),
    .B(_1598_),
    .C(net235),
    .D(_1600_),
    .X(_1866_));
 sky130_fd_sc_hd__and4_1 _5881_ (.A(net260),
    .B(net234),
    .C(_1648_),
    .D(_1796_),
    .X(_1867_));
 sky130_fd_sc_hd__a2111o_1 _5882_ (.A1(\mul_la.lob_4.L[10] ),
    .A2(_1812_),
    .B1(_1865_),
    .C1(_1866_),
    .D1(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__or4_4 _5883_ (.A(_1858_),
    .B(_1863_),
    .C(_1864_),
    .D(_1868_),
    .X(_1869_));
 sky130_fd_sc_hd__and4_1 _5884_ (.A(net264),
    .B(net235),
    .C(_1608_),
    .D(_1789_),
    .X(_1870_));
 sky130_fd_sc_hd__a21o_1 _5885_ (.A1(net262),
    .A2(_1787_),
    .B1(_1870_),
    .X(_1871_));
 sky130_fd_sc_hd__or4_1 _5886_ (.A(_1860_),
    .B(_1865_),
    .C(_1866_),
    .D(_1867_),
    .X(_1872_));
 sky130_fd_sc_hd__o21a_1 _5887_ (.A1(_1871_),
    .A2(_1872_),
    .B1(_1629_),
    .X(_1873_));
 sky130_fd_sc_hd__a21o_1 _5888_ (.A1(\mul_la.lob_4.L[4] ),
    .A2(_1577_),
    .B1(_1859_),
    .X(_1874_));
 sky130_fd_sc_hd__o41a_1 _5889_ (.A1(_1858_),
    .A2(_1861_),
    .A3(_1864_),
    .A4(_1874_),
    .B1(_1629_),
    .X(_1875_));
 sky130_fd_sc_hd__or2_4 _5890_ (.A(_1873_),
    .B(_1875_),
    .X(_1876_));
 sky130_fd_sc_hd__nand2_8 _5891_ (.A(_1629_),
    .B(_1869_),
    .Y(_1877_));
 sky130_fd_sc_hd__or2_1 _5892_ (.A(_1755_),
    .B(_1877_),
    .X(_1878_));
 sky130_fd_sc_hd__nand2_1 _5893_ (.A(net167),
    .B(_1828_),
    .Y(_1879_));
 sky130_fd_sc_hd__and2_1 _5894_ (.A(net257),
    .B(_1703_),
    .X(_1880_));
 sky130_fd_sc_hd__a32o_1 _5895_ (.A1(_1720_),
    .A2(_1758_),
    .A3(_1880_),
    .B1(_1688_),
    .B2(\mul_la.lob_4.L[6] ),
    .X(_1881_));
 sky130_fd_sc_hd__nand2b_2 _5896_ (.A_N(_1702_),
    .B(_1881_),
    .Y(_1882_));
 sky130_fd_sc_hd__a22o_1 _5897_ (.A1(\mul_la.lob_4.L[4] ),
    .A2(_1693_),
    .B1(_1740_),
    .B2(\mul_la.lob_4.L[5] ),
    .X(_1883_));
 sky130_fd_sc_hd__and3_1 _5898_ (.A(net261),
    .B(_1700_),
    .C(_1713_),
    .X(_1884_));
 sky130_fd_sc_hd__a22o_1 _5899_ (.A1(\mul_la.lob_4.L[8] ),
    .A2(_1676_),
    .B1(_1761_),
    .B2(net264),
    .X(_1885_));
 sky130_fd_sc_hd__o21a_1 _5900_ (.A1(_1884_),
    .A2(_1885_),
    .B1(_1704_),
    .X(_1886_));
 sky130_fd_sc_hd__a2111oi_4 _5901_ (.A1(\mul_la.lob_4.L[7] ),
    .A2(_1768_),
    .B1(_1883_),
    .C1(_1886_),
    .D1(_1733_),
    .Y(_1887_));
 sky130_fd_sc_hd__and3_1 _5902_ (.A(net259),
    .B(_1731_),
    .C(_1769_),
    .X(_1888_));
 sky130_fd_sc_hd__a221oi_4 _5903_ (.A1(net263),
    .A2(_1757_),
    .B1(_1773_),
    .B2(net265),
    .C1(_1888_),
    .Y(_1889_));
 sky130_fd_sc_hd__a31oi_4 _5904_ (.A1(_1882_),
    .A2(_1887_),
    .A3(_1889_),
    .B1(_1719_),
    .Y(_1890_));
 sky130_fd_sc_hd__a31o_4 _5905_ (.A1(_1882_),
    .A2(_1887_),
    .A3(_1889_),
    .B1(_1719_),
    .X(_1891_));
 sky130_fd_sc_hd__a2bb2o_1 _5906_ (.A1_N(_1803_),
    .A2_N(net170),
    .B1(_1890_),
    .B2(net188),
    .X(_1892_));
 sky130_fd_sc_hd__and4b_1 _5907_ (.A_N(net171),
    .B(_1890_),
    .C(net188),
    .D(_1804_),
    .X(_1893_));
 sky130_fd_sc_hd__inv_2 _5908_ (.A(_1893_),
    .Y(_1894_));
 sky130_fd_sc_hd__nand2_1 _5909_ (.A(_1892_),
    .B(_1894_),
    .Y(_1895_));
 sky130_fd_sc_hd__xor2_2 _5910_ (.A(_1879_),
    .B(_1895_),
    .X(_1896_));
 sky130_fd_sc_hd__a32o_1 _5911_ (.A1(net167),
    .A2(_1804_),
    .A3(_1848_),
    .B1(_1849_),
    .B2(_1830_),
    .X(_1897_));
 sky130_fd_sc_hd__nand2_1 _5912_ (.A(_1896_),
    .B(_1897_),
    .Y(_1898_));
 sky130_fd_sc_hd__xor2_2 _5913_ (.A(_1896_),
    .B(_1897_),
    .X(_1899_));
 sky130_fd_sc_hd__nand2b_1 _5914_ (.A_N(_1878_),
    .B(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__xnor2_2 _5915_ (.A(_1878_),
    .B(_1899_),
    .Y(_1901_));
 sky130_fd_sc_hd__nand2b_1 _5916_ (.A_N(_1851_),
    .B(_1901_),
    .Y(_1902_));
 sky130_fd_sc_hd__xnor2_1 _5917_ (.A(_1851_),
    .B(_1901_),
    .Y(_1903_));
 sky130_fd_sc_hd__xnor2_1 _5918_ (.A(_1856_),
    .B(_1903_),
    .Y(\mul_la.reg_p[3] ));
 sky130_fd_sc_hd__and4_1 _5919_ (.A(net265),
    .B(_1598_),
    .C(_1599_),
    .D(_1600_),
    .X(_1904_));
 sky130_fd_sc_hd__and4_1 _5920_ (.A(net258),
    .B(_1646_),
    .C(_1648_),
    .D(_1796_),
    .X(_1905_));
 sky130_fd_sc_hd__and4_1 _5921_ (.A(net262),
    .B(_1611_),
    .C(_1617_),
    .D(_1646_),
    .X(_1906_));
 sky130_fd_sc_hd__and4_1 _5922_ (.A(net263),
    .B(net235),
    .C(_1608_),
    .D(_1789_),
    .X(_1907_));
 sky130_fd_sc_hd__or4_1 _5923_ (.A(_1904_),
    .B(_1905_),
    .C(_1906_),
    .D(_1907_),
    .X(_1908_));
 sky130_fd_sc_hd__and2_1 _5924_ (.A(net260),
    .B(_1787_),
    .X(_1909_));
 sky130_fd_sc_hd__and3_1 _5925_ (.A(\mul_la.lob_4.L[8] ),
    .B(_1596_),
    .C(_1611_),
    .X(_1910_));
 sky130_fd_sc_hd__a22o_1 _5926_ (.A1(\mul_la.lob_4.L[5] ),
    .A2(_1577_),
    .B1(_1784_),
    .B2(\mul_la.lob_4.L[6] ),
    .X(_1911_));
 sky130_fd_sc_hd__a32o_1 _5927_ (.A1(net264),
    .A2(_1781_),
    .A3(_1782_),
    .B1(_1818_),
    .B2(\mul_la.lob_4.L[7] ),
    .X(_1912_));
 sky130_fd_sc_hd__a2111o_1 _5928_ (.A1(net255),
    .A2(_1822_),
    .B1(_1910_),
    .C1(_1911_),
    .D1(_1912_),
    .X(_1913_));
 sky130_fd_sc_hd__o31a_4 _5929_ (.A1(_1908_),
    .A2(_1909_),
    .A3(_1913_),
    .B1(_1630_),
    .X(_1914_));
 sky130_fd_sc_hd__inv_2 _5930_ (.A(net186),
    .Y(_1915_));
 sky130_fd_sc_hd__and4b_2 _5931_ (.A_N(_1755_),
    .B(net167),
    .C(_1876_),
    .D(net186),
    .X(_1916_));
 sky130_fd_sc_hd__o22a_1 _5932_ (.A1(_1776_),
    .A2(_1877_),
    .B1(_1915_),
    .B2(_1755_),
    .X(_1917_));
 sky130_fd_sc_hd__nor2_1 _5933_ (.A(_1916_),
    .B(_1917_),
    .Y(_1918_));
 sky130_fd_sc_hd__nor2_1 _5934_ (.A(_1829_),
    .B(net171),
    .Y(_1919_));
 sky130_fd_sc_hd__and4_1 _5935_ (.A(_1686_),
    .B(net233),
    .C(_1703_),
    .D(_1761_),
    .X(_1920_));
 sky130_fd_sc_hd__and3_1 _5936_ (.A(net257),
    .B(_1731_),
    .C(_1769_),
    .X(_1921_));
 sky130_fd_sc_hd__and2_1 _5937_ (.A(net265),
    .B(_1676_),
    .X(_1922_));
 sky130_fd_sc_hd__and4_1 _5938_ (.A(_1686_),
    .B(net233),
    .C(_1703_),
    .D(_1922_),
    .X(_1923_));
 sky130_fd_sc_hd__and2_1 _5939_ (.A(\mul_la.lob_4.L[5] ),
    .B(net232),
    .X(_1924_));
 sky130_fd_sc_hd__and3_1 _5940_ (.A(\mul_la.lob_4.L[6] ),
    .B(_1685_),
    .C(net233),
    .X(_1925_));
 sky130_fd_sc_hd__a2111o_1 _5941_ (.A1(\mul_la.lob_4.L[7] ),
    .A2(_1835_),
    .B1(_1923_),
    .C1(_1924_),
    .D1(_1925_),
    .X(_1926_));
 sky130_fd_sc_hd__and3_1 _5942_ (.A(net259),
    .B(_1700_),
    .C(_1715_),
    .X(_1927_));
 sky130_fd_sc_hd__and3_1 _5943_ (.A(_1672_),
    .B(_1704_),
    .C(_1711_),
    .X(_1928_));
 sky130_fd_sc_hd__and4_1 _5944_ (.A(net263),
    .B(_1672_),
    .C(_1704_),
    .D(_1711_),
    .X(_1929_));
 sky130_fd_sc_hd__a221o_2 _5945_ (.A1(net261),
    .A2(_1757_),
    .B1(_1773_),
    .B2(net264),
    .C1(_1929_),
    .X(_1930_));
 sky130_fd_sc_hd__a32o_1 _5946_ (.A1(\mul_la.lob_4.L[8] ),
    .A2(_1680_),
    .A3(net226),
    .B1(_1758_),
    .B2(_1839_),
    .X(_1931_));
 sky130_fd_sc_hd__or4_4 _5947_ (.A(_1921_),
    .B(_1926_),
    .C(_1927_),
    .D(_1931_),
    .X(_1932_));
 sky130_fd_sc_hd__o21a_4 _5948_ (.A1(_1930_),
    .A2(_1932_),
    .B1(_1720_),
    .X(_1933_));
 sky130_fd_sc_hd__o21ai_4 _5949_ (.A1(_1930_),
    .A2(_1932_),
    .B1(_1720_),
    .Y(_1934_));
 sky130_fd_sc_hd__a22o_1 _5950_ (.A1(_1804_),
    .A2(_1890_),
    .B1(_1933_),
    .B2(net188),
    .X(_1935_));
 sky130_fd_sc_hd__or4_1 _5951_ (.A(_1664_),
    .B(_1803_),
    .C(_1891_),
    .D(net169),
    .X(_1936_));
 sky130_fd_sc_hd__and3_1 _5952_ (.A(_1919_),
    .B(_1935_),
    .C(_1936_),
    .X(_1937_));
 sky130_fd_sc_hd__a21oi_1 _5953_ (.A1(_1935_),
    .A2(_1936_),
    .B1(_1919_),
    .Y(_1938_));
 sky130_fd_sc_hd__a31oi_2 _5954_ (.A1(net167),
    .A2(_1828_),
    .A3(_1892_),
    .B1(_1893_),
    .Y(_1939_));
 sky130_fd_sc_hd__nor3_1 _5955_ (.A(_1937_),
    .B(_1938_),
    .C(_1939_),
    .Y(_1940_));
 sky130_fd_sc_hd__or3_1 _5956_ (.A(_1937_),
    .B(_1938_),
    .C(_1939_),
    .X(_1941_));
 sky130_fd_sc_hd__o21ai_1 _5957_ (.A1(_1937_),
    .A2(_1938_),
    .B1(_1939_),
    .Y(_1942_));
 sky130_fd_sc_hd__and3_1 _5958_ (.A(_1918_),
    .B(_1941_),
    .C(_1942_),
    .X(_1943_));
 sky130_fd_sc_hd__a21oi_1 _5959_ (.A1(_1941_),
    .A2(_1942_),
    .B1(_1918_),
    .Y(_1944_));
 sky130_fd_sc_hd__or2_1 _5960_ (.A(_1943_),
    .B(_1944_),
    .X(_1945_));
 sky130_fd_sc_hd__a21o_1 _5961_ (.A1(_1898_),
    .A2(_1900_),
    .B1(_1945_),
    .X(_1946_));
 sky130_fd_sc_hd__nand3_1 _5962_ (.A(_1898_),
    .B(_1900_),
    .C(_1945_),
    .Y(_1947_));
 sky130_fd_sc_hd__nand2_1 _5963_ (.A(_1946_),
    .B(_1947_),
    .Y(_1948_));
 sky130_fd_sc_hd__or2_1 _5964_ (.A(_1902_),
    .B(_1948_),
    .X(_1949_));
 sky130_fd_sc_hd__nand2_1 _5965_ (.A(_1902_),
    .B(_1948_),
    .Y(_1950_));
 sky130_fd_sc_hd__nand2_1 _5966_ (.A(_1949_),
    .B(_1950_),
    .Y(_1951_));
 sky130_fd_sc_hd__nor2_1 _5967_ (.A(_1855_),
    .B(_1901_),
    .Y(_1952_));
 sky130_fd_sc_hd__or2_1 _5968_ (.A(_1951_),
    .B(_1952_),
    .X(_1953_));
 sky130_fd_sc_hd__nand2_1 _5969_ (.A(_1948_),
    .B(_1952_),
    .Y(_1954_));
 sky130_fd_sc_hd__and2_1 _5970_ (.A(net251),
    .B(_1954_),
    .X(_1955_));
 sky130_fd_sc_hd__a2bb2o_1 _5971_ (.A1_N(net251),
    .A2_N(_1951_),
    .B1(_1953_),
    .B2(_1955_),
    .X(\mul_la.reg_p[4] ));
 sky130_fd_sc_hd__a211o_1 _5972_ (.A1(_1766_),
    .A2(_1774_),
    .B1(_1915_),
    .C1(_1725_),
    .X(_1956_));
 sky130_fd_sc_hd__nor2_1 _5973_ (.A(net171),
    .B(_1877_),
    .Y(_1957_));
 sky130_fd_sc_hd__xnor2_1 _5974_ (.A(_1956_),
    .B(_1957_),
    .Y(_1958_));
 sky130_fd_sc_hd__a22o_1 _5975_ (.A1(net264),
    .A2(_1779_),
    .B1(_1812_),
    .B2(net262),
    .X(_1959_));
 sky130_fd_sc_hd__a22o_1 _5976_ (.A1(\mul_la.lob_4.L[6] ),
    .A2(net236),
    .B1(_1784_),
    .B2(\mul_la.lob_4.L[7] ),
    .X(_1960_));
 sky130_fd_sc_hd__and2_1 _5977_ (.A(net258),
    .B(_1787_),
    .X(_1961_));
 sky130_fd_sc_hd__and3_1 _5978_ (.A(net263),
    .B(_1781_),
    .C(_1782_),
    .X(_1962_));
 sky130_fd_sc_hd__and4_1 _5979_ (.A(net255),
    .B(_1610_),
    .C(net234),
    .D(_1648_),
    .X(_1963_));
 sky130_fd_sc_hd__a211o_1 _5980_ (.A1(net260),
    .A2(_1777_),
    .B1(_1960_),
    .C1(_1963_),
    .X(_1964_));
 sky130_fd_sc_hd__a221o_1 _5981_ (.A1(net265),
    .A2(_1798_),
    .B1(_1818_),
    .B2(\mul_la.lob_4.L[8] ),
    .C1(_1962_),
    .X(_1965_));
 sky130_fd_sc_hd__o41a_4 _5982_ (.A1(_1959_),
    .A2(_1961_),
    .A3(_1964_),
    .A4(_1965_),
    .B1(_1625_),
    .X(_1966_));
 sky130_fd_sc_hd__o41ai_4 _5983_ (.A1(_1959_),
    .A2(_1961_),
    .A3(_1964_),
    .A4(_1965_),
    .B1(_1625_),
    .Y(_1967_));
 sky130_fd_sc_hd__nor2_1 _5984_ (.A(_1755_),
    .B(_1967_),
    .Y(_1968_));
 sky130_fd_sc_hd__xor2_1 _5985_ (.A(_1958_),
    .B(_1968_),
    .X(_1969_));
 sky130_fd_sc_hd__nor2_1 _5986_ (.A(_1829_),
    .B(_1891_),
    .Y(_1970_));
 sky130_fd_sc_hd__a32o_1 _5987_ (.A1(net265),
    .A2(_1680_),
    .A3(_1689_),
    .B1(_1685_),
    .B2(\mul_la.lob_4.L[7] ),
    .X(_1971_));
 sky130_fd_sc_hd__a32o_1 _5988_ (.A1(net256),
    .A2(_1695_),
    .A3(_1731_),
    .B1(\mul_la.lob_4.L[6] ),
    .B2(net232),
    .X(_1972_));
 sky130_fd_sc_hd__a22o_1 _5989_ (.A1(net264),
    .A2(_1676_),
    .B1(_1761_),
    .B2(net261),
    .X(_1973_));
 sky130_fd_sc_hd__a22o_1 _5990_ (.A1(\mul_la.lob_4.L[8] ),
    .A2(_1835_),
    .B1(_1973_),
    .B2(_1704_),
    .X(_1974_));
 sky130_fd_sc_hd__a211o_2 _5991_ (.A1(_1695_),
    .A2(_1971_),
    .B1(_1972_),
    .C1(_1974_),
    .X(_1975_));
 sky130_fd_sc_hd__and3_1 _5992_ (.A(net257),
    .B(_1700_),
    .C(_1715_),
    .X(_1976_));
 sky130_fd_sc_hd__a221o_4 _5993_ (.A1(net259),
    .A2(_1757_),
    .B1(_1773_),
    .B2(net263),
    .C1(_1976_),
    .X(_1977_));
 sky130_fd_sc_hd__o21a_2 _5994_ (.A1(_1975_),
    .A2(_1977_),
    .B1(_1709_),
    .X(_1978_));
 sky130_fd_sc_hd__o21ai_2 _5995_ (.A1(_1975_),
    .A2(_1977_),
    .B1(_1709_),
    .Y(_1979_));
 sky130_fd_sc_hd__a22o_1 _5996_ (.A1(_1804_),
    .A2(_1933_),
    .B1(_1978_),
    .B2(net187),
    .X(_1980_));
 sky130_fd_sc_hd__or4_1 _5997_ (.A(_1664_),
    .B(_1803_),
    .C(net169),
    .D(net168),
    .X(_1981_));
 sky130_fd_sc_hd__nand3_1 _5998_ (.A(_1970_),
    .B(_1980_),
    .C(_1981_),
    .Y(_1982_));
 sky130_fd_sc_hd__a21o_1 _5999_ (.A1(_1980_),
    .A2(_1981_),
    .B1(_1970_),
    .X(_1983_));
 sky130_fd_sc_hd__a21bo_1 _6000_ (.A1(_1919_),
    .A2(_1935_),
    .B1_N(_1936_),
    .X(_1984_));
 sky130_fd_sc_hd__nand3_2 _6001_ (.A(_1982_),
    .B(_1983_),
    .C(_1984_),
    .Y(_1985_));
 sky130_fd_sc_hd__a21o_1 _6002_ (.A1(_1982_),
    .A2(_1983_),
    .B1(_1984_),
    .X(_1986_));
 sky130_fd_sc_hd__nand3_2 _6003_ (.A(_1969_),
    .B(_1985_),
    .C(_1986_),
    .Y(_1987_));
 sky130_fd_sc_hd__a21o_1 _6004_ (.A1(_1985_),
    .A2(_1986_),
    .B1(_1969_),
    .X(_1988_));
 sky130_fd_sc_hd__o211a_1 _6005_ (.A1(_1940_),
    .A2(_1943_),
    .B1(_1987_),
    .C1(_1988_),
    .X(_1989_));
 sky130_fd_sc_hd__a211o_1 _6006_ (.A1(_1987_),
    .A2(_1988_),
    .B1(_1940_),
    .C1(_1943_),
    .X(_1990_));
 sky130_fd_sc_hd__and2b_1 _6007_ (.A_N(_1989_),
    .B(_1990_),
    .X(_1991_));
 sky130_fd_sc_hd__xnor2_2 _6008_ (.A(_1916_),
    .B(_1991_),
    .Y(_1992_));
 sky130_fd_sc_hd__nand2_1 _6009_ (.A(_1946_),
    .B(_1949_),
    .Y(_1993_));
 sky130_fd_sc_hd__xnor2_1 _6010_ (.A(_1992_),
    .B(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__xor2_1 _6011_ (.A(_1955_),
    .B(_1994_),
    .X(\mul_la.reg_p[5] ));
 sky130_fd_sc_hd__a21o_1 _6012_ (.A1(_1916_),
    .A2(_1990_),
    .B1(_1989_),
    .X(_1995_));
 sky130_fd_sc_hd__a32o_1 _6013_ (.A1(net167),
    .A2(net186),
    .A3(_1957_),
    .B1(_1958_),
    .B2(_1968_),
    .X(_1996_));
 sky130_fd_sc_hd__and3_1 _6014_ (.A(net262),
    .B(_1781_),
    .C(_1782_),
    .X(_1997_));
 sky130_fd_sc_hd__a22o_1 _6015_ (.A1(\mul_la.lob_4.L[7] ),
    .A2(net236),
    .B1(_1784_),
    .B2(\mul_la.lob_4.L[8] ),
    .X(_1998_));
 sky130_fd_sc_hd__and3_1 _6016_ (.A(\mul_la.lob_4.L[10] ),
    .B(_1596_),
    .C(_1611_),
    .X(_1999_));
 sky130_fd_sc_hd__and2_1 _6017_ (.A(net265),
    .B(_1818_),
    .X(_2000_));
 sky130_fd_sc_hd__and4_1 _6018_ (.A(net255),
    .B(_1598_),
    .C(net235),
    .D(_1619_),
    .X(_2001_));
 sky130_fd_sc_hd__and4_1 _6019_ (.A(net258),
    .B(_1611_),
    .C(_1617_),
    .D(net234),
    .X(_2002_));
 sky130_fd_sc_hd__a2111o_2 _6020_ (.A1(\mul_la.lob_4.L[11] ),
    .A2(_1779_),
    .B1(_1997_),
    .C1(_1999_),
    .D1(_2001_),
    .X(_2003_));
 sky130_fd_sc_hd__a2111o_2 _6021_ (.A1(net260),
    .A2(_1812_),
    .B1(_1998_),
    .C1(_2000_),
    .D1(_2002_),
    .X(_2004_));
 sky130_fd_sc_hd__o21a_4 _6022_ (.A1(_2003_),
    .A2(_2004_),
    .B1(_1621_),
    .X(_2005_));
 sky130_fd_sc_hd__o21ai_4 _6023_ (.A1(_2003_),
    .A2(_2004_),
    .B1(_1621_),
    .Y(_2006_));
 sky130_fd_sc_hd__nor2_1 _6024_ (.A(_1755_),
    .B(_2006_),
    .Y(_2007_));
 sky130_fd_sc_hd__nand2_1 _6025_ (.A(_1996_),
    .B(_2007_),
    .Y(_2008_));
 sky130_fd_sc_hd__xor2_1 _6026_ (.A(_1996_),
    .B(_2007_),
    .X(_2009_));
 sky130_fd_sc_hd__nor2_1 _6027_ (.A(net171),
    .B(_1915_),
    .Y(_2010_));
 sky130_fd_sc_hd__nor2_1 _6028_ (.A(_1877_),
    .B(_1891_),
    .Y(_2011_));
 sky130_fd_sc_hd__xnor2_1 _6029_ (.A(_2010_),
    .B(_2011_),
    .Y(_2012_));
 sky130_fd_sc_hd__nand2_1 _6030_ (.A(_1775_),
    .B(_1966_),
    .Y(_2013_));
 sky130_fd_sc_hd__or2_1 _6031_ (.A(_2012_),
    .B(_2013_),
    .X(_2014_));
 sky130_fd_sc_hd__xor2_1 _6032_ (.A(_2012_),
    .B(_2013_),
    .X(_2015_));
 sky130_fd_sc_hd__nor2_1 _6033_ (.A(_1829_),
    .B(net169),
    .Y(_2016_));
 sky130_fd_sc_hd__a32o_1 _6034_ (.A1(net263),
    .A2(_1676_),
    .A3(_1703_),
    .B1(_1688_),
    .B2(net265),
    .X(_2017_));
 sky130_fd_sc_hd__and4b_1 _6035_ (.A_N(_1688_),
    .B(_1680_),
    .C(net264),
    .D(_1686_),
    .X(_2018_));
 sky130_fd_sc_hd__and2_1 _6036_ (.A(\mul_la.lob_4.L[8] ),
    .B(_1685_),
    .X(_2019_));
 sky130_fd_sc_hd__a211o_1 _6037_ (.A1(_1686_),
    .A2(_2017_),
    .B1(_2018_),
    .C1(_2019_),
    .X(_2020_));
 sky130_fd_sc_hd__a22o_1 _6038_ (.A1(\mul_la.lob_4.L[7] ),
    .A2(net232),
    .B1(_1715_),
    .B2(net256),
    .X(_2021_));
 sky130_fd_sc_hd__a221o_4 _6039_ (.A1(net257),
    .A2(_1757_),
    .B1(_1928_),
    .B2(net259),
    .C1(_2021_),
    .X(_2022_));
 sky130_fd_sc_hd__a22o_4 _6040_ (.A1(net261),
    .A2(_1773_),
    .B1(_2020_),
    .B2(net233),
    .X(_2023_));
 sky130_fd_sc_hd__o21a_4 _6041_ (.A1(_2022_),
    .A2(_2023_),
    .B1(_1700_),
    .X(_2024_));
 sky130_fd_sc_hd__o21ai_4 _6042_ (.A1(_2022_),
    .A2(_2023_),
    .B1(_1700_),
    .Y(_2025_));
 sky130_fd_sc_hd__a22o_1 _6043_ (.A1(_1804_),
    .A2(_1978_),
    .B1(_2024_),
    .B2(net187),
    .X(_2026_));
 sky130_fd_sc_hd__or4_1 _6044_ (.A(_1664_),
    .B(_1803_),
    .C(net168),
    .D(_2025_),
    .X(_2027_));
 sky130_fd_sc_hd__nand3_1 _6045_ (.A(_2016_),
    .B(_2026_),
    .C(_2027_),
    .Y(_2028_));
 sky130_fd_sc_hd__a21o_1 _6046_ (.A1(_2026_),
    .A2(_2027_),
    .B1(_2016_),
    .X(_2029_));
 sky130_fd_sc_hd__a21bo_1 _6047_ (.A1(_1970_),
    .A2(_1980_),
    .B1_N(_1981_),
    .X(_2030_));
 sky130_fd_sc_hd__and3_1 _6048_ (.A(_2028_),
    .B(_2029_),
    .C(_2030_),
    .X(_2031_));
 sky130_fd_sc_hd__nand3_1 _6049_ (.A(_2028_),
    .B(_2029_),
    .C(_2030_),
    .Y(_2032_));
 sky130_fd_sc_hd__a21o_1 _6050_ (.A1(_2028_),
    .A2(_2029_),
    .B1(_2030_),
    .X(_2033_));
 sky130_fd_sc_hd__and3_1 _6051_ (.A(_2015_),
    .B(_2032_),
    .C(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__a21oi_1 _6052_ (.A1(_2032_),
    .A2(_2033_),
    .B1(_2015_),
    .Y(_2035_));
 sky130_fd_sc_hd__a211o_1 _6053_ (.A1(_1985_),
    .A2(_1987_),
    .B1(_2034_),
    .C1(_2035_),
    .X(_2036_));
 sky130_fd_sc_hd__o211ai_1 _6054_ (.A1(_2034_),
    .A2(_2035_),
    .B1(_1985_),
    .C1(_1987_),
    .Y(_2037_));
 sky130_fd_sc_hd__nand3_1 _6055_ (.A(_2009_),
    .B(_2036_),
    .C(_2037_),
    .Y(_2038_));
 sky130_fd_sc_hd__a21o_1 _6056_ (.A1(_2036_),
    .A2(_2037_),
    .B1(_2009_),
    .X(_2039_));
 sky130_fd_sc_hd__and3_1 _6057_ (.A(_1995_),
    .B(_2038_),
    .C(_2039_),
    .X(_2040_));
 sky130_fd_sc_hd__a21oi_1 _6058_ (.A1(_2038_),
    .A2(_2039_),
    .B1(_1995_),
    .Y(_2041_));
 sky130_fd_sc_hd__nor4_2 _6059_ (.A(_1946_),
    .B(_1992_),
    .C(_2040_),
    .D(_2041_),
    .Y(_2042_));
 sky130_fd_sc_hd__inv_2 _6060_ (.A(net166),
    .Y(_2043_));
 sky130_fd_sc_hd__o22a_1 _6061_ (.A1(_1946_),
    .A2(_1992_),
    .B1(_2040_),
    .B2(_2041_),
    .X(_2044_));
 sky130_fd_sc_hd__nor2_1 _6062_ (.A(_2042_),
    .B(_2044_),
    .Y(_2045_));
 sky130_fd_sc_hd__nor2_1 _6063_ (.A(_1949_),
    .B(_1992_),
    .Y(_2046_));
 sky130_fd_sc_hd__or3b_1 _6064_ (.A(_1949_),
    .B(_1992_),
    .C_N(_2045_),
    .X(_2047_));
 sky130_fd_sc_hd__xnor2_1 _6065_ (.A(_2045_),
    .B(_2046_),
    .Y(_2048_));
 sky130_fd_sc_hd__o21a_1 _6066_ (.A1(_1954_),
    .A2(_1994_),
    .B1(net251),
    .X(_2049_));
 sky130_fd_sc_hd__xnor2_1 _6067_ (.A(_2048_),
    .B(_2049_),
    .Y(\mul_la.reg_p[6] ));
 sky130_fd_sc_hd__or3b_2 _6068_ (.A(_1954_),
    .B(_1994_),
    .C_N(_2048_),
    .X(_2050_));
 sky130_fd_sc_hd__nand2_1 _6069_ (.A(net700),
    .B(_2050_),
    .Y(_2051_));
 sky130_fd_sc_hd__a21bo_1 _6070_ (.A1(_2010_),
    .A2(_2011_),
    .B1_N(_2014_),
    .X(_2052_));
 sky130_fd_sc_hd__and2_2 _6071_ (.A(net255),
    .B(_1611_),
    .X(_2053_));
 sky130_fd_sc_hd__a32o_1 _6072_ (.A1(net263),
    .A2(_1596_),
    .A3(_1611_),
    .B1(_1818_),
    .B2(\mul_la.lob_4.L[10] ),
    .X(_2054_));
 sky130_fd_sc_hd__a21oi_2 _6073_ (.A1(net234),
    .A2(_2053_),
    .B1(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__and4_1 _6074_ (.A(net262),
    .B(_1598_),
    .C(net235),
    .D(_1600_),
    .X(_2056_));
 sky130_fd_sc_hd__and4_1 _6075_ (.A(net258),
    .B(net235),
    .C(_1608_),
    .D(_1789_),
    .X(_2057_));
 sky130_fd_sc_hd__and3_1 _6076_ (.A(net259),
    .B(_1781_),
    .C(_1782_),
    .X(_2058_));
 sky130_fd_sc_hd__a22o_1 _6077_ (.A1(\mul_la.lob_4.L[8] ),
    .A2(net236),
    .B1(_1784_),
    .B2(\mul_la.lob_4.L[9] ),
    .X(_2059_));
 sky130_fd_sc_hd__nor4_1 _6078_ (.A(_2056_),
    .B(_2057_),
    .C(_2058_),
    .D(_2059_),
    .Y(_2060_));
 sky130_fd_sc_hd__a21oi_4 _6079_ (.A1(_2055_),
    .A2(net215),
    .B1(_1618_),
    .Y(_2061_));
 sky130_fd_sc_hd__a21o_4 _6080_ (.A1(_2055_),
    .A2(_2060_),
    .B1(_1618_),
    .X(_2062_));
 sky130_fd_sc_hd__nor2_1 _6081_ (.A(_1755_),
    .B(_2062_),
    .Y(_2063_));
 sky130_fd_sc_hd__and3_1 _6082_ (.A(_1775_),
    .B(_2005_),
    .C(_2063_),
    .X(_2064_));
 sky130_fd_sc_hd__a21o_1 _6083_ (.A1(_1775_),
    .A2(_2005_),
    .B1(_2063_),
    .X(_2065_));
 sky130_fd_sc_hd__and2b_1 _6084_ (.A_N(_2064_),
    .B(_2065_),
    .X(_2066_));
 sky130_fd_sc_hd__and2_1 _6085_ (.A(_2052_),
    .B(_2066_),
    .X(_2067_));
 sky130_fd_sc_hd__xnor2_1 _6086_ (.A(_2052_),
    .B(_2066_),
    .Y(_2068_));
 sky130_fd_sc_hd__nor2_1 _6087_ (.A(net170),
    .B(net184),
    .Y(_2069_));
 sky130_fd_sc_hd__a22o_1 _6088_ (.A1(_1890_),
    .A2(net186),
    .B1(_1933_),
    .B2(_1876_),
    .X(_2070_));
 sky130_fd_sc_hd__or4_1 _6089_ (.A(_1877_),
    .B(_1891_),
    .C(_1915_),
    .D(net169),
    .X(_2071_));
 sky130_fd_sc_hd__nand2_1 _6090_ (.A(_2070_),
    .B(_2071_),
    .Y(_2072_));
 sky130_fd_sc_hd__xnor2_1 _6091_ (.A(_2069_),
    .B(_2072_),
    .Y(_2073_));
 sky130_fd_sc_hd__nor2_1 _6092_ (.A(_1829_),
    .B(net168),
    .Y(_2074_));
 sky130_fd_sc_hd__and4_1 _6093_ (.A(net259),
    .B(_1670_),
    .C(_1681_),
    .D(_1696_),
    .X(_2075_));
 sky130_fd_sc_hd__nand2_1 _6094_ (.A(net264),
    .B(_1688_),
    .Y(_2076_));
 sky130_fd_sc_hd__a2111o_1 _6095_ (.A1(_1678_),
    .A2(_1679_),
    .B1(_1688_),
    .C1(_1675_),
    .D1(_3374_),
    .X(_2077_));
 sky130_fd_sc_hd__a211oi_1 _6096_ (.A1(_2076_),
    .A2(_2077_),
    .B1(_1685_),
    .C1(net232),
    .Y(_2078_));
 sky130_fd_sc_hd__a22o_1 _6097_ (.A1(\mul_la.lob_4.L[8] ),
    .A2(net232),
    .B1(_1694_),
    .B2(\mul_la.lob_4.L[7] ),
    .X(_2079_));
 sky130_fd_sc_hd__a211o_1 _6098_ (.A1(net257),
    .A2(_1920_),
    .B1(_2078_),
    .C1(_2079_),
    .X(_2080_));
 sky130_fd_sc_hd__and2_1 _6099_ (.A(net265),
    .B(_1685_),
    .X(_2081_));
 sky130_fd_sc_hd__and4b_1 _6100_ (.A_N(_1688_),
    .B(_1680_),
    .C(net263),
    .D(_1686_),
    .X(_2082_));
 sky130_fd_sc_hd__o21a_1 _6101_ (.A1(_2081_),
    .A2(_2082_),
    .B1(_1695_),
    .X(_2083_));
 sky130_fd_sc_hd__and3_1 _6102_ (.A(net256),
    .B(_1696_),
    .C(_1727_),
    .X(_2084_));
 sky130_fd_sc_hd__o41a_2 _6103_ (.A1(_2075_),
    .A2(_2080_),
    .A3(_2083_),
    .A4(_2084_),
    .B1(_1699_),
    .X(_2085_));
 sky130_fd_sc_hd__a22o_1 _6104_ (.A1(_1804_),
    .A2(_2024_),
    .B1(net182),
    .B2(net187),
    .X(_2086_));
 sky130_fd_sc_hd__or4b_1 _6105_ (.A(_1664_),
    .B(_1803_),
    .C(_2025_),
    .D_N(net182),
    .X(_2087_));
 sky130_fd_sc_hd__nand3_1 _6106_ (.A(_2074_),
    .B(_2086_),
    .C(_2087_),
    .Y(_2088_));
 sky130_fd_sc_hd__a21o_1 _6107_ (.A1(_2086_),
    .A2(_2087_),
    .B1(_2074_),
    .X(_2089_));
 sky130_fd_sc_hd__a21bo_1 _6108_ (.A1(_2016_),
    .A2(_2026_),
    .B1_N(_2027_),
    .X(_2090_));
 sky130_fd_sc_hd__nand3_1 _6109_ (.A(_2088_),
    .B(_2089_),
    .C(_2090_),
    .Y(_2091_));
 sky130_fd_sc_hd__a21o_1 _6110_ (.A1(_2088_),
    .A2(_2089_),
    .B1(_2090_),
    .X(_2092_));
 sky130_fd_sc_hd__nand3_1 _6111_ (.A(_2073_),
    .B(_2091_),
    .C(_2092_),
    .Y(_2093_));
 sky130_fd_sc_hd__a21o_1 _6112_ (.A1(_2091_),
    .A2(_2092_),
    .B1(_2073_),
    .X(_2094_));
 sky130_fd_sc_hd__o211a_1 _6113_ (.A1(_2031_),
    .A2(_2034_),
    .B1(_2093_),
    .C1(_2094_),
    .X(_2095_));
 sky130_fd_sc_hd__a211oi_2 _6114_ (.A1(_2093_),
    .A2(_2094_),
    .B1(_2031_),
    .C1(_2034_),
    .Y(_2096_));
 sky130_fd_sc_hd__nor3_1 _6115_ (.A(_2068_),
    .B(_2095_),
    .C(_2096_),
    .Y(_2097_));
 sky130_fd_sc_hd__o21a_1 _6116_ (.A1(_2095_),
    .A2(_2096_),
    .B1(_2068_),
    .X(_2098_));
 sky130_fd_sc_hd__a211oi_1 _6117_ (.A1(_2036_),
    .A2(_2038_),
    .B1(_2097_),
    .C1(_2098_),
    .Y(_2099_));
 sky130_fd_sc_hd__o211a_1 _6118_ (.A1(_2097_),
    .A2(_2098_),
    .B1(_2036_),
    .C1(_2038_),
    .X(_2100_));
 sky130_fd_sc_hd__or3_1 _6119_ (.A(_2008_),
    .B(_2099_),
    .C(_2100_),
    .X(_2101_));
 sky130_fd_sc_hd__o21ai_1 _6120_ (.A1(_2099_),
    .A2(_2100_),
    .B1(_2008_),
    .Y(_2102_));
 sky130_fd_sc_hd__nand2_1 _6121_ (.A(_2101_),
    .B(_2102_),
    .Y(_2103_));
 sky130_fd_sc_hd__nor2_1 _6122_ (.A(_2040_),
    .B(net166),
    .Y(_2104_));
 sky130_fd_sc_hd__xnor2_1 _6123_ (.A(_2103_),
    .B(_2104_),
    .Y(_2105_));
 sky130_fd_sc_hd__nor2_1 _6124_ (.A(_2047_),
    .B(_2105_),
    .Y(_2106_));
 sky130_fd_sc_hd__and2_1 _6125_ (.A(_2047_),
    .B(_2105_),
    .X(_2107_));
 sky130_fd_sc_hd__nor2_1 _6126_ (.A(_2106_),
    .B(_2107_),
    .Y(_2108_));
 sky130_fd_sc_hd__xnor2_1 _6127_ (.A(_2051_),
    .B(_2108_),
    .Y(\mul_la.reg_p[7] ));
 sky130_fd_sc_hd__and3_1 _6128_ (.A(_2040_),
    .B(_2101_),
    .C(_2102_),
    .X(_2109_));
 sky130_fd_sc_hd__a21bo_1 _6129_ (.A1(_2069_),
    .A2(_2070_),
    .B1_N(_2071_),
    .X(_2110_));
 sky130_fd_sc_hd__and3_1 _6130_ (.A(net258),
    .B(_1781_),
    .C(_1782_),
    .X(_2111_));
 sky130_fd_sc_hd__a32o_1 _6131_ (.A1(net255),
    .A2(net235),
    .A3(_1789_),
    .B1(_1818_),
    .B2(\mul_la.lob_4.L[11] ),
    .X(_2112_));
 sky130_fd_sc_hd__a22o_1 _6132_ (.A1(\mul_la.lob_4.L[9] ),
    .A2(net236),
    .B1(_1784_),
    .B2(\mul_la.lob_4.L[10] ),
    .X(_2113_));
 sky130_fd_sc_hd__a221o_1 _6133_ (.A1(net260),
    .A2(_1779_),
    .B1(_1798_),
    .B2(net262),
    .C1(_2113_),
    .X(_2114_));
 sky130_fd_sc_hd__o31ai_4 _6134_ (.A1(_2111_),
    .A2(_2112_),
    .A3(_2114_),
    .B1(_1608_),
    .Y(_2115_));
 sky130_fd_sc_hd__inv_2 _6135_ (.A(_2115_),
    .Y(_2116_));
 sky130_fd_sc_hd__nor2_1 _6136_ (.A(_1755_),
    .B(net181),
    .Y(_2117_));
 sky130_fd_sc_hd__a211o_1 _6137_ (.A1(_1766_),
    .A2(_1774_),
    .B1(_2062_),
    .C1(_1725_),
    .X(_2118_));
 sky130_fd_sc_hd__nor2_1 _6138_ (.A(net171),
    .B(_2006_),
    .Y(_2119_));
 sky130_fd_sc_hd__xnor2_2 _6139_ (.A(_2118_),
    .B(_2119_),
    .Y(_2120_));
 sky130_fd_sc_hd__xnor2_2 _6140_ (.A(_2117_),
    .B(_2120_),
    .Y(_2121_));
 sky130_fd_sc_hd__and2b_1 _6141_ (.A_N(_2121_),
    .B(_2110_),
    .X(_2122_));
 sky130_fd_sc_hd__xnor2_2 _6142_ (.A(_2110_),
    .B(_2121_),
    .Y(_2123_));
 sky130_fd_sc_hd__and2_1 _6143_ (.A(_2064_),
    .B(_2123_),
    .X(_2124_));
 sky130_fd_sc_hd__xnor2_2 _6144_ (.A(_2064_),
    .B(_2123_),
    .Y(_2125_));
 sky130_fd_sc_hd__nand2_2 _6145_ (.A(_1890_),
    .B(_1966_),
    .Y(_2126_));
 sky130_fd_sc_hd__a22o_1 _6146_ (.A1(net186),
    .A2(_1933_),
    .B1(_1978_),
    .B2(_1876_),
    .X(_2127_));
 sky130_fd_sc_hd__or4_1 _6147_ (.A(_1877_),
    .B(_1915_),
    .C(_1934_),
    .D(net168),
    .X(_2128_));
 sky130_fd_sc_hd__nand2_1 _6148_ (.A(_2127_),
    .B(_2128_),
    .Y(_2129_));
 sky130_fd_sc_hd__xor2_2 _6149_ (.A(_2126_),
    .B(_2129_),
    .X(_2130_));
 sky130_fd_sc_hd__nand2_1 _6150_ (.A(_1828_),
    .B(_2024_),
    .Y(_2131_));
 sky130_fd_sc_hd__a21boi_2 _6151_ (.A1(_1794_),
    .A2(_1802_),
    .B1_N(net183),
    .Y(_2132_));
 sky130_fd_sc_hd__and4_2 _6152_ (.A(net257),
    .B(_1670_),
    .C(_1681_),
    .D(net226),
    .X(_2133_));
 sky130_fd_sc_hd__and3_2 _6153_ (.A(net261),
    .B(_1680_),
    .C(net226),
    .X(_2134_));
 sky130_fd_sc_hd__nor2_1 _6154_ (.A(_3373_),
    .B(_1675_),
    .Y(_2135_));
 sky130_fd_sc_hd__and3b_1 _6155_ (.A_N(_1670_),
    .B(_1675_),
    .C(net256),
    .X(_2136_));
 sky130_fd_sc_hd__o2111a_1 _6156_ (.A1(_2135_),
    .A2(_2136_),
    .B1(_1686_),
    .C1(net233),
    .D1(_1703_),
    .X(_2137_));
 sky130_fd_sc_hd__and2_1 _6157_ (.A(net265),
    .B(net232),
    .X(_2138_));
 sky130_fd_sc_hd__and3_1 _6158_ (.A(net264),
    .B(_1685_),
    .C(net233),
    .X(_2139_));
 sky130_fd_sc_hd__a2111o_2 _6159_ (.A1(net263),
    .A2(_1835_),
    .B1(_2137_),
    .C1(_2138_),
    .D1(_2139_),
    .X(_2140_));
 sky130_fd_sc_hd__o31a_4 _6160_ (.A1(_2133_),
    .A2(_2134_),
    .A3(_2140_),
    .B1(_1672_),
    .X(_2141_));
 sky130_fd_sc_hd__o31ai_4 _6161_ (.A1(_2133_),
    .A2(_2134_),
    .A3(_2140_),
    .B1(_1672_),
    .Y(_2142_));
 sky130_fd_sc_hd__nand2_1 _6162_ (.A(net187),
    .B(_2141_),
    .Y(_2143_));
 sky130_fd_sc_hd__and3_1 _6163_ (.A(net187),
    .B(_2132_),
    .C(_2141_),
    .X(_2144_));
 sky130_fd_sc_hd__xnor2_2 _6164_ (.A(_2132_),
    .B(_2143_),
    .Y(_2145_));
 sky130_fd_sc_hd__xnor2_2 _6165_ (.A(_2131_),
    .B(_2145_),
    .Y(_2146_));
 sky130_fd_sc_hd__a21boi_2 _6166_ (.A1(_2074_),
    .A2(_2086_),
    .B1_N(_2087_),
    .Y(_2147_));
 sky130_fd_sc_hd__nand2b_1 _6167_ (.A_N(_2147_),
    .B(_2146_),
    .Y(_2148_));
 sky130_fd_sc_hd__xnor2_2 _6168_ (.A(_2146_),
    .B(_2147_),
    .Y(_2149_));
 sky130_fd_sc_hd__xnor2_2 _6169_ (.A(_2130_),
    .B(_2149_),
    .Y(_2150_));
 sky130_fd_sc_hd__a21bo_1 _6170_ (.A1(_2073_),
    .A2(_2092_),
    .B1_N(_2091_),
    .X(_2151_));
 sky130_fd_sc_hd__nand2b_1 _6171_ (.A_N(_2150_),
    .B(_2151_),
    .Y(_2152_));
 sky130_fd_sc_hd__xor2_2 _6172_ (.A(_2150_),
    .B(_2151_),
    .X(_2153_));
 sky130_fd_sc_hd__xor2_2 _6173_ (.A(_2125_),
    .B(_2153_),
    .X(_2154_));
 sky130_fd_sc_hd__o21ba_1 _6174_ (.A1(_2068_),
    .A2(_2096_),
    .B1_N(_2095_),
    .X(_2155_));
 sky130_fd_sc_hd__and2b_1 _6175_ (.A_N(_2155_),
    .B(_2154_),
    .X(_2156_));
 sky130_fd_sc_hd__xnor2_2 _6176_ (.A(_2154_),
    .B(_2155_),
    .Y(_2157_));
 sky130_fd_sc_hd__xor2_2 _6177_ (.A(_2067_),
    .B(_2157_),
    .X(_2158_));
 sky130_fd_sc_hd__o21ba_1 _6178_ (.A1(_2008_),
    .A2(_2100_),
    .B1_N(_2099_),
    .X(_2159_));
 sky130_fd_sc_hd__nand2b_1 _6179_ (.A_N(_2159_),
    .B(_2158_),
    .Y(_2160_));
 sky130_fd_sc_hd__xnor2_2 _6180_ (.A(_2158_),
    .B(_2159_),
    .Y(_2161_));
 sky130_fd_sc_hd__nand2_1 _6181_ (.A(_2109_),
    .B(_2161_),
    .Y(_2162_));
 sky130_fd_sc_hd__xnor2_2 _6182_ (.A(_2109_),
    .B(_2161_),
    .Y(_2163_));
 sky130_fd_sc_hd__nor2_1 _6183_ (.A(_2043_),
    .B(_2103_),
    .Y(_2164_));
 sky130_fd_sc_hd__or3_1 _6184_ (.A(_2043_),
    .B(_2103_),
    .C(_2163_),
    .X(_2165_));
 sky130_fd_sc_hd__xnor2_2 _6185_ (.A(_2163_),
    .B(_2164_),
    .Y(_2166_));
 sky130_fd_sc_hd__xnor2_1 _6186_ (.A(_2106_),
    .B(_2166_),
    .Y(_2167_));
 sky130_fd_sc_hd__o21a_1 _6187_ (.A1(_2050_),
    .A2(_2108_),
    .B1(net700),
    .X(_2168_));
 sky130_fd_sc_hd__xnor2_1 _6188_ (.A(_2167_),
    .B(_2168_),
    .Y(\mul_la.reg_p[8] ));
 sky130_fd_sc_hd__or3b_1 _6189_ (.A(_2050_),
    .B(_2108_),
    .C_N(_2167_),
    .X(_2169_));
 sky130_fd_sc_hd__nand2_1 _6190_ (.A(net251),
    .B(_2169_),
    .Y(_2170_));
 sky130_fd_sc_hd__and4_1 _6191_ (.A(net258),
    .B(_1598_),
    .C(_1599_),
    .D(_1600_),
    .X(_2171_));
 sky130_fd_sc_hd__a32o_1 _6192_ (.A1(net260),
    .A2(_1596_),
    .A3(_1611_),
    .B1(_1818_),
    .B2(net262),
    .X(_2172_));
 sky130_fd_sc_hd__a22o_1 _6193_ (.A1(\mul_la.lob_4.L[10] ),
    .A2(net236),
    .B1(_1784_),
    .B2(\mul_la.lob_4.L[11] ),
    .X(_2173_));
 sky130_fd_sc_hd__and3_1 _6194_ (.A(net256),
    .B(_1610_),
    .C(_1781_),
    .X(_2174_));
 sky130_fd_sc_hd__o41a_4 _6195_ (.A1(_2171_),
    .A2(_2172_),
    .A3(_2173_),
    .A4(_2174_),
    .B1(_1604_),
    .X(_2175_));
 sky130_fd_sc_hd__inv_2 _6196_ (.A(net214),
    .Y(_2176_));
 sky130_fd_sc_hd__nor2_1 _6197_ (.A(_1755_),
    .B(_2176_),
    .Y(_2177_));
 sky130_fd_sc_hd__o21a_1 _6198_ (.A1(_2122_),
    .A2(_2124_),
    .B1(_2177_),
    .X(_2178_));
 sky130_fd_sc_hd__nor3_1 _6199_ (.A(_2122_),
    .B(_2124_),
    .C(_2177_),
    .Y(_2179_));
 sky130_fd_sc_hd__nor2_1 _6200_ (.A(_2178_),
    .B(_2179_),
    .Y(_2180_));
 sky130_fd_sc_hd__a32o_1 _6201_ (.A1(_1775_),
    .A2(_2061_),
    .A3(_2119_),
    .B1(_2120_),
    .B2(_2117_),
    .X(_2181_));
 sky130_fd_sc_hd__o21ai_2 _6202_ (.A1(_2126_),
    .A2(_2129_),
    .B1(_2128_),
    .Y(_2182_));
 sky130_fd_sc_hd__nor2_1 _6203_ (.A(_1776_),
    .B(net181),
    .Y(_2183_));
 sky130_fd_sc_hd__or2_1 _6204_ (.A(net170),
    .B(_2062_),
    .X(_2184_));
 sky130_fd_sc_hd__nand2_2 _6205_ (.A(_1890_),
    .B(_2005_),
    .Y(_2185_));
 sky130_fd_sc_hd__xnor2_2 _6206_ (.A(_2184_),
    .B(_2185_),
    .Y(_2186_));
 sky130_fd_sc_hd__or3_1 _6207_ (.A(_1776_),
    .B(net181),
    .C(_2186_),
    .X(_2187_));
 sky130_fd_sc_hd__xnor2_2 _6208_ (.A(_2183_),
    .B(_2186_),
    .Y(_2188_));
 sky130_fd_sc_hd__and2_1 _6209_ (.A(_2182_),
    .B(_2188_),
    .X(_2189_));
 sky130_fd_sc_hd__xnor2_2 _6210_ (.A(_2182_),
    .B(_2188_),
    .Y(_2190_));
 sky130_fd_sc_hd__and2b_1 _6211_ (.A_N(_2190_),
    .B(_2181_),
    .X(_2191_));
 sky130_fd_sc_hd__xnor2_2 _6212_ (.A(_2181_),
    .B(_2190_),
    .Y(_2192_));
 sky130_fd_sc_hd__nor2_1 _6213_ (.A(net169),
    .B(net184),
    .Y(_2193_));
 sky130_fd_sc_hd__a22o_1 _6214_ (.A1(net186),
    .A2(_1978_),
    .B1(_2024_),
    .B2(_1876_),
    .X(_2194_));
 sky130_fd_sc_hd__or4_1 _6215_ (.A(_1877_),
    .B(_1915_),
    .C(_1979_),
    .D(_2025_),
    .X(_2195_));
 sky130_fd_sc_hd__nand2_1 _6216_ (.A(_2194_),
    .B(_2195_),
    .Y(_2196_));
 sky130_fd_sc_hd__xor2_2 _6217_ (.A(_2193_),
    .B(_2196_),
    .X(_2197_));
 sky130_fd_sc_hd__nand2_1 _6218_ (.A(net172),
    .B(net182),
    .Y(_2198_));
 sky130_fd_sc_hd__a21oi_2 _6219_ (.A1(_1794_),
    .A2(_1802_),
    .B1(net180),
    .Y(_2199_));
 sky130_fd_sc_hd__a22o_1 _6220_ (.A1(net259),
    .A2(_1680_),
    .B1(_1681_),
    .B2(net256),
    .X(_2200_));
 sky130_fd_sc_hd__a22o_2 _6221_ (.A1(net264),
    .A2(net232),
    .B1(_1740_),
    .B2(\mul_la.lob_4.L[11] ),
    .X(_2201_));
 sky130_fd_sc_hd__a32o_1 _6222_ (.A1(net257),
    .A2(_1676_),
    .A3(_1703_),
    .B1(_1688_),
    .B2(net261),
    .X(_2202_));
 sky130_fd_sc_hd__a32o_2 _6223_ (.A1(_1686_),
    .A2(net233),
    .A3(_2202_),
    .B1(_2200_),
    .B2(net226),
    .X(_2203_));
 sky130_fd_sc_hd__o21a_4 _6224_ (.A1(_2201_),
    .A2(_2203_),
    .B1(_1670_),
    .X(_2204_));
 sky130_fd_sc_hd__o21ai_4 _6225_ (.A1(_2201_),
    .A2(_2203_),
    .B1(_1670_),
    .Y(_2205_));
 sky130_fd_sc_hd__nand2_1 _6226_ (.A(net187),
    .B(_2204_),
    .Y(_2206_));
 sky130_fd_sc_hd__and3_1 _6227_ (.A(net187),
    .B(_2199_),
    .C(_2204_),
    .X(_2207_));
 sky130_fd_sc_hd__xnor2_2 _6228_ (.A(_2199_),
    .B(_2206_),
    .Y(_2208_));
 sky130_fd_sc_hd__xnor2_2 _6229_ (.A(_2198_),
    .B(_2208_),
    .Y(_2209_));
 sky130_fd_sc_hd__a31o_1 _6230_ (.A1(net172),
    .A2(_2024_),
    .A3(_2145_),
    .B1(_2144_),
    .X(_2210_));
 sky130_fd_sc_hd__nand2_1 _6231_ (.A(_2209_),
    .B(_2210_),
    .Y(_2211_));
 sky130_fd_sc_hd__nor2_1 _6232_ (.A(_2209_),
    .B(_2210_),
    .Y(_2212_));
 sky130_fd_sc_hd__xor2_1 _6233_ (.A(_2209_),
    .B(_2210_),
    .X(_2213_));
 sky130_fd_sc_hd__xnor2_2 _6234_ (.A(_2197_),
    .B(_2213_),
    .Y(_2214_));
 sky130_fd_sc_hd__a21bo_1 _6235_ (.A1(_2130_),
    .A2(_2149_),
    .B1_N(_2148_),
    .X(_2215_));
 sky130_fd_sc_hd__nand2_1 _6236_ (.A(_2214_),
    .B(_2215_),
    .Y(_2216_));
 sky130_fd_sc_hd__xor2_2 _6237_ (.A(_2214_),
    .B(_2215_),
    .X(_2217_));
 sky130_fd_sc_hd__xor2_2 _6238_ (.A(_2192_),
    .B(_2217_),
    .X(_2218_));
 sky130_fd_sc_hd__o21a_1 _6239_ (.A1(_2125_),
    .A2(_2153_),
    .B1(_2152_),
    .X(_2219_));
 sky130_fd_sc_hd__and2b_1 _6240_ (.A_N(_2219_),
    .B(_2218_),
    .X(_2220_));
 sky130_fd_sc_hd__xnor2_2 _6241_ (.A(_2218_),
    .B(_2219_),
    .Y(_2221_));
 sky130_fd_sc_hd__xnor2_2 _6242_ (.A(_2180_),
    .B(_2221_),
    .Y(_2222_));
 sky130_fd_sc_hd__a21oi_2 _6243_ (.A1(_2067_),
    .A2(_2157_),
    .B1(_2156_),
    .Y(_2223_));
 sky130_fd_sc_hd__nor2_1 _6244_ (.A(_2222_),
    .B(_2223_),
    .Y(_2224_));
 sky130_fd_sc_hd__xnor2_2 _6245_ (.A(_2222_),
    .B(_2223_),
    .Y(_2225_));
 sky130_fd_sc_hd__a21boi_1 _6246_ (.A1(_2109_),
    .A2(_2161_),
    .B1_N(_2160_),
    .Y(_2226_));
 sky130_fd_sc_hd__xnor2_2 _6247_ (.A(_2225_),
    .B(_2226_),
    .Y(_2227_));
 sky130_fd_sc_hd__a21boi_1 _6248_ (.A1(_2106_),
    .A2(_2166_),
    .B1_N(_2165_),
    .Y(_2228_));
 sky130_fd_sc_hd__xor2_1 _6249_ (.A(_2227_),
    .B(_2228_),
    .X(_2229_));
 sky130_fd_sc_hd__xnor2_1 _6250_ (.A(_2170_),
    .B(_2229_),
    .Y(\mul_la.reg_p[9] ));
 sky130_fd_sc_hd__nand2_1 _6251_ (.A(net167),
    .B(net214),
    .Y(_2230_));
 sky130_fd_sc_hd__a22o_1 _6252_ (.A1(\mul_la.lob_4.L[11] ),
    .A2(net236),
    .B1(_1784_),
    .B2(net261),
    .X(_2231_));
 sky130_fd_sc_hd__and3_1 _6253_ (.A(net256),
    .B(_1598_),
    .C(net235),
    .X(_2232_));
 sky130_fd_sc_hd__a32o_1 _6254_ (.A1(net258),
    .A2(_1596_),
    .A3(_1611_),
    .B1(_1818_),
    .B2(net260),
    .X(_2233_));
 sky130_fd_sc_hd__o31a_4 _6255_ (.A1(_2231_),
    .A2(_2232_),
    .A3(_2233_),
    .B1(_1600_),
    .X(_2234_));
 sky130_fd_sc_hd__inv_2 _6256_ (.A(net213),
    .Y(_2235_));
 sky130_fd_sc_hd__or2_1 _6257_ (.A(_1755_),
    .B(_2235_),
    .X(_2236_));
 sky130_fd_sc_hd__nor2_2 _6258_ (.A(_2230_),
    .B(_2236_),
    .Y(_2237_));
 sky130_fd_sc_hd__xor2_1 _6259_ (.A(_2230_),
    .B(_2236_),
    .X(_2238_));
 sky130_fd_sc_hd__o21a_2 _6260_ (.A1(_2189_),
    .A2(_2191_),
    .B1(_2238_),
    .X(_2239_));
 sky130_fd_sc_hd__nor3_1 _6261_ (.A(_2189_),
    .B(_2191_),
    .C(_2238_),
    .Y(_2240_));
 sky130_fd_sc_hd__nor2_1 _6262_ (.A(_2239_),
    .B(_2240_),
    .Y(_2241_));
 sky130_fd_sc_hd__o31ai_4 _6263_ (.A1(net171),
    .A2(_2062_),
    .A3(_2185_),
    .B1(_2187_),
    .Y(_2242_));
 sky130_fd_sc_hd__a21bo_1 _6264_ (.A1(_2193_),
    .A2(_2194_),
    .B1_N(_2195_),
    .X(_2243_));
 sky130_fd_sc_hd__nand2_1 _6265_ (.A(_1890_),
    .B(_2061_),
    .Y(_2244_));
 sky130_fd_sc_hd__nor2_1 _6266_ (.A(net169),
    .B(_2006_),
    .Y(_2245_));
 sky130_fd_sc_hd__xnor2_2 _6267_ (.A(_2244_),
    .B(_2245_),
    .Y(_2246_));
 sky130_fd_sc_hd__nor2_1 _6268_ (.A(net170),
    .B(net181),
    .Y(_2247_));
 sky130_fd_sc_hd__xnor2_2 _6269_ (.A(_2246_),
    .B(_2247_),
    .Y(_2248_));
 sky130_fd_sc_hd__and2b_1 _6270_ (.A_N(_2248_),
    .B(_2243_),
    .X(_2249_));
 sky130_fd_sc_hd__xnor2_2 _6271_ (.A(_2243_),
    .B(_2248_),
    .Y(_2250_));
 sky130_fd_sc_hd__xor2_2 _6272_ (.A(_2242_),
    .B(_2250_),
    .X(_2251_));
 sky130_fd_sc_hd__nor2_1 _6273_ (.A(net184),
    .B(net168),
    .Y(_2252_));
 sky130_fd_sc_hd__a22o_1 _6274_ (.A1(net186),
    .A2(_2024_),
    .B1(net183),
    .B2(_1876_),
    .X(_2253_));
 sky130_fd_sc_hd__or4b_1 _6275_ (.A(_1877_),
    .B(_1915_),
    .C(_2025_),
    .D_N(net182),
    .X(_2254_));
 sky130_fd_sc_hd__and3_1 _6276_ (.A(_2252_),
    .B(_2253_),
    .C(_2254_),
    .X(_2255_));
 sky130_fd_sc_hd__a21oi_1 _6277_ (.A1(_2253_),
    .A2(_2254_),
    .B1(_2252_),
    .Y(_2256_));
 sky130_fd_sc_hd__or2_2 _6278_ (.A(_2255_),
    .B(_2256_),
    .X(_2257_));
 sky130_fd_sc_hd__nand2_1 _6279_ (.A(net172),
    .B(_2141_),
    .Y(_2258_));
 sky130_fd_sc_hd__a21oi_2 _6280_ (.A1(_1794_),
    .A2(_1802_),
    .B1(_2205_),
    .Y(_2259_));
 sky130_fd_sc_hd__and3_2 _6281_ (.A(net257),
    .B(_1680_),
    .C(net226),
    .X(_2260_));
 sky130_fd_sc_hd__and2_1 _6282_ (.A(net263),
    .B(net232),
    .X(_2261_));
 sky130_fd_sc_hd__and3_1 _6283_ (.A(net261),
    .B(_1685_),
    .C(net233),
    .X(_2262_));
 sky130_fd_sc_hd__a2111o_2 _6284_ (.A1(net259),
    .A2(_1835_),
    .B1(_1839_),
    .C1(_2261_),
    .D1(_2262_),
    .X(_2263_));
 sky130_fd_sc_hd__o21a_4 _6285_ (.A1(_2260_),
    .A2(_2263_),
    .B1(_1676_),
    .X(_2264_));
 sky130_fd_sc_hd__o21ai_4 _6286_ (.A1(_2260_),
    .A2(_2263_),
    .B1(_1676_),
    .Y(_2265_));
 sky130_fd_sc_hd__nand2_1 _6287_ (.A(net187),
    .B(_2264_),
    .Y(_2266_));
 sky130_fd_sc_hd__and3_1 _6288_ (.A(net187),
    .B(_2259_),
    .C(_2264_),
    .X(_2267_));
 sky130_fd_sc_hd__xnor2_2 _6289_ (.A(_2259_),
    .B(_2266_),
    .Y(_2268_));
 sky130_fd_sc_hd__xnor2_2 _6290_ (.A(_2258_),
    .B(_2268_),
    .Y(_2269_));
 sky130_fd_sc_hd__a31o_1 _6291_ (.A1(net172),
    .A2(net182),
    .A3(_2208_),
    .B1(_2207_),
    .X(_2270_));
 sky130_fd_sc_hd__nand2_1 _6292_ (.A(_2269_),
    .B(_2270_),
    .Y(_2271_));
 sky130_fd_sc_hd__nor2_1 _6293_ (.A(_2269_),
    .B(_2270_),
    .Y(_2272_));
 sky130_fd_sc_hd__xor2_1 _6294_ (.A(_2269_),
    .B(_2270_),
    .X(_2273_));
 sky130_fd_sc_hd__xnor2_2 _6295_ (.A(_2257_),
    .B(_2273_),
    .Y(_2274_));
 sky130_fd_sc_hd__o21a_1 _6296_ (.A1(_2197_),
    .A2(_2212_),
    .B1(_2211_),
    .X(_2275_));
 sky130_fd_sc_hd__nand2b_1 _6297_ (.A_N(_2275_),
    .B(_2274_),
    .Y(_2276_));
 sky130_fd_sc_hd__xnor2_2 _6298_ (.A(_2274_),
    .B(_2275_),
    .Y(_2277_));
 sky130_fd_sc_hd__xnor2_2 _6299_ (.A(_2251_),
    .B(_2277_),
    .Y(_2278_));
 sky130_fd_sc_hd__a21bo_1 _6300_ (.A1(_2192_),
    .A2(_2217_),
    .B1_N(_2216_),
    .X(_2279_));
 sky130_fd_sc_hd__and2b_1 _6301_ (.A_N(_2278_),
    .B(_2279_),
    .X(_2280_));
 sky130_fd_sc_hd__xnor2_2 _6302_ (.A(_2278_),
    .B(_2279_),
    .Y(_2281_));
 sky130_fd_sc_hd__xnor2_2 _6303_ (.A(_2241_),
    .B(_2281_),
    .Y(_2282_));
 sky130_fd_sc_hd__a21oi_2 _6304_ (.A1(_2180_),
    .A2(_2221_),
    .B1(_2220_),
    .Y(_2283_));
 sky130_fd_sc_hd__nor2_1 _6305_ (.A(_2282_),
    .B(_2283_),
    .Y(_2284_));
 sky130_fd_sc_hd__xor2_2 _6306_ (.A(_2282_),
    .B(_2283_),
    .X(_2285_));
 sky130_fd_sc_hd__xor2_2 _6307_ (.A(_2178_),
    .B(_2285_),
    .X(_2286_));
 sky130_fd_sc_hd__nor2_1 _6308_ (.A(_2160_),
    .B(_2225_),
    .Y(_2287_));
 sky130_fd_sc_hd__or2_1 _6309_ (.A(_2224_),
    .B(_2287_),
    .X(_2288_));
 sky130_fd_sc_hd__xnor2_1 _6310_ (.A(_2286_),
    .B(_2288_),
    .Y(_2289_));
 sky130_fd_sc_hd__or4b_2 _6311_ (.A(_2047_),
    .B(_2105_),
    .C(_2227_),
    .D_N(_2166_),
    .X(_2290_));
 sky130_fd_sc_hd__o22a_1 _6312_ (.A1(_2162_),
    .A2(_2225_),
    .B1(_2227_),
    .B2(_2165_),
    .X(_2291_));
 sky130_fd_sc_hd__nand3_1 _6313_ (.A(_2289_),
    .B(_2290_),
    .C(_2291_),
    .Y(_2292_));
 sky130_fd_sc_hd__a21o_1 _6314_ (.A1(_2290_),
    .A2(_2291_),
    .B1(_2289_),
    .X(_2293_));
 sky130_fd_sc_hd__nand2_1 _6315_ (.A(_2292_),
    .B(_2293_),
    .Y(_2294_));
 sky130_fd_sc_hd__nor2_1 _6316_ (.A(_2169_),
    .B(_2229_),
    .Y(_2295_));
 sky130_fd_sc_hd__nor2_1 _6317_ (.A(_1809_),
    .B(_2295_),
    .Y(_2296_));
 sky130_fd_sc_hd__xnor2_1 _6318_ (.A(_2294_),
    .B(_2296_),
    .Y(\mul_la.reg_p[10] ));
 sky130_fd_sc_hd__a21oi_1 _6319_ (.A1(_2294_),
    .A2(_2295_),
    .B1(_1809_),
    .Y(_2297_));
 sky130_fd_sc_hd__nand2_1 _6320_ (.A(_2286_),
    .B(_2287_),
    .Y(_2298_));
 sky130_fd_sc_hd__a21oi_2 _6321_ (.A1(_2242_),
    .A2(_2250_),
    .B1(_2249_),
    .Y(_2299_));
 sky130_fd_sc_hd__a32o_1 _6322_ (.A1(net260),
    .A2(_1584_),
    .A3(_1610_),
    .B1(net262),
    .B2(net236),
    .X(_2300_));
 sky130_fd_sc_hd__a31o_1 _6323_ (.A1(net258),
    .A2(_1586_),
    .A3(_1641_),
    .B1(_2300_),
    .X(_2301_));
 sky130_fd_sc_hd__o21a_4 _6324_ (.A1(_2053_),
    .A2(_2301_),
    .B1(_1596_),
    .X(_2302_));
 sky130_fd_sc_hd__o21ai_4 _6325_ (.A1(_2053_),
    .A2(_2301_),
    .B1(_1596_),
    .Y(_2303_));
 sky130_fd_sc_hd__nor2_1 _6326_ (.A(_1755_),
    .B(net179),
    .Y(_2304_));
 sky130_fd_sc_hd__nor2_1 _6327_ (.A(net170),
    .B(_2176_),
    .Y(_2305_));
 sky130_fd_sc_hd__a21oi_1 _6328_ (.A1(net167),
    .A2(_2234_),
    .B1(_2305_),
    .Y(_2306_));
 sky130_fd_sc_hd__a21o_1 _6329_ (.A1(net167),
    .A2(_2234_),
    .B1(_2305_),
    .X(_2307_));
 sky130_fd_sc_hd__and3_1 _6330_ (.A(net167),
    .B(_2234_),
    .C(_2305_),
    .X(_2308_));
 sky130_fd_sc_hd__nor2_1 _6331_ (.A(_2306_),
    .B(_2308_),
    .Y(_2309_));
 sky130_fd_sc_hd__xnor2_2 _6332_ (.A(_2304_),
    .B(_2309_),
    .Y(_2310_));
 sky130_fd_sc_hd__inv_2 _6333_ (.A(_2310_),
    .Y(_2311_));
 sky130_fd_sc_hd__nand2_1 _6334_ (.A(_2237_),
    .B(_2311_),
    .Y(_2312_));
 sky130_fd_sc_hd__xor2_2 _6335_ (.A(_2237_),
    .B(_2310_),
    .X(_2313_));
 sky130_fd_sc_hd__nor2_1 _6336_ (.A(_2299_),
    .B(_2313_),
    .Y(_2314_));
 sky130_fd_sc_hd__xor2_2 _6337_ (.A(_2299_),
    .B(_2313_),
    .X(_2315_));
 sky130_fd_sc_hd__a32o_1 _6338_ (.A1(_1890_),
    .A2(_2061_),
    .A3(_2245_),
    .B1(_2246_),
    .B2(_2247_),
    .X(_2316_));
 sky130_fd_sc_hd__a21bo_1 _6339_ (.A1(_2252_),
    .A2(_2253_),
    .B1_N(_2254_),
    .X(_2317_));
 sky130_fd_sc_hd__nor2_1 _6340_ (.A(_1891_),
    .B(net181),
    .Y(_2318_));
 sky130_fd_sc_hd__nor2_2 _6341_ (.A(net169),
    .B(_2062_),
    .Y(_2319_));
 sky130_fd_sc_hd__nor2_2 _6342_ (.A(net168),
    .B(_2006_),
    .Y(_2320_));
 sky130_fd_sc_hd__nand2_1 _6343_ (.A(_2319_),
    .B(_2320_),
    .Y(_2321_));
 sky130_fd_sc_hd__xnor2_4 _6344_ (.A(_2319_),
    .B(_2320_),
    .Y(_2322_));
 sky130_fd_sc_hd__xnor2_2 _6345_ (.A(_2318_),
    .B(_2322_),
    .Y(_2323_));
 sky130_fd_sc_hd__and2_1 _6346_ (.A(_2317_),
    .B(_2323_),
    .X(_2324_));
 sky130_fd_sc_hd__xor2_2 _6347_ (.A(_2317_),
    .B(_2323_),
    .X(_2325_));
 sky130_fd_sc_hd__xor2_2 _6348_ (.A(_2316_),
    .B(_2325_),
    .X(_2326_));
 sky130_fd_sc_hd__nor2_1 _6349_ (.A(net184),
    .B(_2025_),
    .Y(_2327_));
 sky130_fd_sc_hd__nand2_1 _6350_ (.A(net186),
    .B(net182),
    .Y(_2328_));
 sky130_fd_sc_hd__nor2_1 _6351_ (.A(_1877_),
    .B(net180),
    .Y(_2329_));
 sky130_fd_sc_hd__and3_1 _6352_ (.A(_1914_),
    .B(net183),
    .C(_2329_),
    .X(_2330_));
 sky130_fd_sc_hd__xnor2_2 _6353_ (.A(_2328_),
    .B(_2329_),
    .Y(_2331_));
 sky130_fd_sc_hd__xor2_2 _6354_ (.A(_2327_),
    .B(_2331_),
    .X(_2332_));
 sky130_fd_sc_hd__nand2_1 _6355_ (.A(net172),
    .B(_2204_),
    .Y(_2333_));
 sky130_fd_sc_hd__a21oi_2 _6356_ (.A1(_1794_),
    .A2(_1802_),
    .B1(_2265_),
    .Y(_2334_));
 sky130_fd_sc_hd__and2_2 _6357_ (.A(net257),
    .B(_1835_),
    .X(_2335_));
 sky130_fd_sc_hd__nor2_1 _6358_ (.A(_3374_),
    .B(_1692_),
    .Y(_2336_));
 sky130_fd_sc_hd__a221o_2 _6359_ (.A1(net256),
    .A2(net226),
    .B1(_1740_),
    .B2(net259),
    .C1(_2336_),
    .X(_2337_));
 sky130_fd_sc_hd__o21a_4 _6360_ (.A1(_2335_),
    .A2(_2337_),
    .B1(_1680_),
    .X(_2338_));
 sky130_fd_sc_hd__o21ai_4 _6361_ (.A1(_2335_),
    .A2(_2337_),
    .B1(_1680_),
    .Y(_2339_));
 sky130_fd_sc_hd__nand2_1 _6362_ (.A(net187),
    .B(_2338_),
    .Y(_2340_));
 sky130_fd_sc_hd__and3_1 _6363_ (.A(net187),
    .B(_2334_),
    .C(_2338_),
    .X(_2341_));
 sky130_fd_sc_hd__xnor2_2 _6364_ (.A(_2334_),
    .B(_2340_),
    .Y(_2342_));
 sky130_fd_sc_hd__xnor2_2 _6365_ (.A(_2333_),
    .B(_2342_),
    .Y(_2343_));
 sky130_fd_sc_hd__a31o_1 _6366_ (.A1(net172),
    .A2(_2141_),
    .A3(_2268_),
    .B1(_2267_),
    .X(_2344_));
 sky130_fd_sc_hd__and2_1 _6367_ (.A(_2343_),
    .B(_2344_),
    .X(_2345_));
 sky130_fd_sc_hd__xor2_2 _6368_ (.A(_2343_),
    .B(_2344_),
    .X(_2346_));
 sky130_fd_sc_hd__xnor2_2 _6369_ (.A(_2332_),
    .B(_2346_),
    .Y(_2347_));
 sky130_fd_sc_hd__o21ai_2 _6370_ (.A1(_2257_),
    .A2(_2272_),
    .B1(_2271_),
    .Y(_2348_));
 sky130_fd_sc_hd__nand2b_1 _6371_ (.A_N(_2347_),
    .B(_2348_),
    .Y(_2349_));
 sky130_fd_sc_hd__xnor2_2 _6372_ (.A(_2347_),
    .B(_2348_),
    .Y(_2350_));
 sky130_fd_sc_hd__xnor2_2 _6373_ (.A(_2326_),
    .B(_2350_),
    .Y(_2351_));
 sky130_fd_sc_hd__a21bo_1 _6374_ (.A1(_2251_),
    .A2(_2277_),
    .B1_N(_2276_),
    .X(_2352_));
 sky130_fd_sc_hd__and2b_1 _6375_ (.A_N(_2351_),
    .B(_2352_),
    .X(_2353_));
 sky130_fd_sc_hd__xnor2_2 _6376_ (.A(_2351_),
    .B(_2352_),
    .Y(_2354_));
 sky130_fd_sc_hd__xnor2_2 _6377_ (.A(_2315_),
    .B(_2354_),
    .Y(_2355_));
 sky130_fd_sc_hd__a21oi_2 _6378_ (.A1(_2241_),
    .A2(_2281_),
    .B1(_2280_),
    .Y(_2356_));
 sky130_fd_sc_hd__nor2_1 _6379_ (.A(_2355_),
    .B(_2356_),
    .Y(_2357_));
 sky130_fd_sc_hd__xor2_2 _6380_ (.A(_2355_),
    .B(_2356_),
    .X(_2358_));
 sky130_fd_sc_hd__xor2_2 _6381_ (.A(_2239_),
    .B(_2358_),
    .X(_2359_));
 sky130_fd_sc_hd__a21oi_2 _6382_ (.A1(_2178_),
    .A2(_2285_),
    .B1(_2284_),
    .Y(_2360_));
 sky130_fd_sc_hd__nand2b_1 _6383_ (.A_N(_2360_),
    .B(_2359_),
    .Y(_2361_));
 sky130_fd_sc_hd__xnor2_2 _6384_ (.A(_2359_),
    .B(_2360_),
    .Y(_2362_));
 sky130_fd_sc_hd__inv_2 _6385_ (.A(_2362_),
    .Y(_2363_));
 sky130_fd_sc_hd__and3_1 _6386_ (.A(_2224_),
    .B(_2286_),
    .C(_2362_),
    .X(_2364_));
 sky130_fd_sc_hd__nand3_1 _6387_ (.A(_2224_),
    .B(_2286_),
    .C(_2362_),
    .Y(_2365_));
 sky130_fd_sc_hd__a21oi_1 _6388_ (.A1(_2224_),
    .A2(_2286_),
    .B1(_2362_),
    .Y(_2366_));
 sky130_fd_sc_hd__or2_1 _6389_ (.A(_2364_),
    .B(_2366_),
    .X(_2367_));
 sky130_fd_sc_hd__and3_1 _6390_ (.A(_2293_),
    .B(_2298_),
    .C(_2367_),
    .X(_2368_));
 sky130_fd_sc_hd__a21oi_1 _6391_ (.A1(_2293_),
    .A2(_2298_),
    .B1(_2367_),
    .Y(_2369_));
 sky130_fd_sc_hd__or2_1 _6392_ (.A(_2368_),
    .B(_2369_),
    .X(_2370_));
 sky130_fd_sc_hd__xnor2_1 _6393_ (.A(_2297_),
    .B(_2370_),
    .Y(\mul_la.reg_p[11] ));
 sky130_fd_sc_hd__a21oi_2 _6394_ (.A1(_2239_),
    .A2(_2358_),
    .B1(_2357_),
    .Y(_2371_));
 sky130_fd_sc_hd__a21o_2 _6395_ (.A1(_2316_),
    .A2(_2325_),
    .B1(_2324_),
    .X(_2372_));
 sky130_fd_sc_hd__nand2_1 _6396_ (.A(net255),
    .B(_1641_),
    .Y(_2373_));
 sky130_fd_sc_hd__nand2_1 _6397_ (.A(net260),
    .B(net236),
    .Y(_2374_));
 sky130_fd_sc_hd__nand2_1 _6398_ (.A(net258),
    .B(_1784_),
    .Y(_2375_));
 sky130_fd_sc_hd__a31oi_4 _6399_ (.A1(_2373_),
    .A2(_2374_),
    .A3(_2375_),
    .B1(_1587_),
    .Y(_2376_));
 sky130_fd_sc_hd__a31o_1 _6400_ (.A1(_2373_),
    .A2(_2374_),
    .A3(_2375_),
    .B1(_1587_),
    .X(_2377_));
 sky130_fd_sc_hd__or2_2 _6401_ (.A(_1755_),
    .B(net178),
    .X(_2378_));
 sky130_fd_sc_hd__nand2_2 _6402_ (.A(net167),
    .B(_2302_),
    .Y(_2379_));
 sky130_fd_sc_hd__o22a_1 _6403_ (.A1(_1891_),
    .A2(_2176_),
    .B1(_2235_),
    .B2(net170),
    .X(_2380_));
 sky130_fd_sc_hd__and4b_1 _6404_ (.A_N(net170),
    .B(_1890_),
    .C(_2175_),
    .D(_2234_),
    .X(_2381_));
 sky130_fd_sc_hd__nor2_2 _6405_ (.A(_2380_),
    .B(_2381_),
    .Y(_2382_));
 sky130_fd_sc_hd__xnor2_4 _6406_ (.A(_2379_),
    .B(_2382_),
    .Y(_2383_));
 sky130_fd_sc_hd__a21o_1 _6407_ (.A1(_2304_),
    .A2(_2307_),
    .B1(_2308_),
    .X(_2384_));
 sky130_fd_sc_hd__and2_1 _6408_ (.A(_2383_),
    .B(_2384_),
    .X(_2385_));
 sky130_fd_sc_hd__xor2_4 _6409_ (.A(_2383_),
    .B(_2384_),
    .X(_2386_));
 sky130_fd_sc_hd__xnor2_4 _6410_ (.A(_2378_),
    .B(_2386_),
    .Y(_2387_));
 sky130_fd_sc_hd__xor2_4 _6411_ (.A(_2372_),
    .B(_2387_),
    .X(_2388_));
 sky130_fd_sc_hd__xnor2_2 _6412_ (.A(_2312_),
    .B(_2388_),
    .Y(_2389_));
 sky130_fd_sc_hd__o31ai_4 _6413_ (.A1(_1891_),
    .A2(net181),
    .A3(_2322_),
    .B1(_2321_),
    .Y(_2390_));
 sky130_fd_sc_hd__a21oi_2 _6414_ (.A1(_2327_),
    .A2(_2331_),
    .B1(_2330_),
    .Y(_2391_));
 sky130_fd_sc_hd__o22a_1 _6415_ (.A1(_2006_),
    .A2(_2025_),
    .B1(_2062_),
    .B2(net168),
    .X(_2392_));
 sky130_fd_sc_hd__or4_2 _6416_ (.A(net168),
    .B(_2006_),
    .C(_2025_),
    .D(_2062_),
    .X(_2393_));
 sky130_fd_sc_hd__nand2b_1 _6417_ (.A_N(_2392_),
    .B(_2393_),
    .Y(_2394_));
 sky130_fd_sc_hd__nor2_1 _6418_ (.A(net169),
    .B(net181),
    .Y(_2395_));
 sky130_fd_sc_hd__xnor2_2 _6419_ (.A(_2394_),
    .B(_2395_),
    .Y(_2396_));
 sky130_fd_sc_hd__nand2b_1 _6420_ (.A_N(_2391_),
    .B(_2396_),
    .Y(_2397_));
 sky130_fd_sc_hd__xnor2_2 _6421_ (.A(_2391_),
    .B(_2396_),
    .Y(_2398_));
 sky130_fd_sc_hd__xnor2_2 _6422_ (.A(_2390_),
    .B(_2398_),
    .Y(_2399_));
 sky130_fd_sc_hd__nand2_1 _6423_ (.A(_1914_),
    .B(_2141_),
    .Y(_2400_));
 sky130_fd_sc_hd__and3_1 _6424_ (.A(_1629_),
    .B(_1869_),
    .C(_2204_),
    .X(_2401_));
 sky130_fd_sc_hd__and3_1 _6425_ (.A(_1914_),
    .B(_2141_),
    .C(_2401_),
    .X(_2402_));
 sky130_fd_sc_hd__xnor2_1 _6426_ (.A(_2400_),
    .B(_2401_),
    .Y(_2403_));
 sky130_fd_sc_hd__and3_1 _6427_ (.A(_1966_),
    .B(net183),
    .C(_2403_),
    .X(_2404_));
 sky130_fd_sc_hd__a21oi_1 _6428_ (.A1(_1966_),
    .A2(net183),
    .B1(_2403_),
    .Y(_2405_));
 sky130_fd_sc_hd__nor2_1 _6429_ (.A(_2404_),
    .B(_2405_),
    .Y(_2406_));
 sky130_fd_sc_hd__nand2_1 _6430_ (.A(net172),
    .B(_2264_),
    .Y(_2407_));
 sky130_fd_sc_hd__a21oi_2 _6431_ (.A1(_1794_),
    .A2(_1802_),
    .B1(_2339_),
    .Y(_2408_));
 sky130_fd_sc_hd__o21a_1 _6432_ (.A1(net259),
    .A2(net233),
    .B1(_1688_),
    .X(_2409_));
 sky130_fd_sc_hd__o221a_4 _6433_ (.A1(net256),
    .A2(_1702_),
    .B1(_1741_),
    .B2(net257),
    .C1(_2409_),
    .X(_2410_));
 sky130_fd_sc_hd__o221ai_4 _6434_ (.A1(net256),
    .A2(_1702_),
    .B1(_1741_),
    .B2(net257),
    .C1(_2409_),
    .Y(_2411_));
 sky130_fd_sc_hd__nand2_1 _6435_ (.A(net188),
    .B(_2410_),
    .Y(_2412_));
 sky130_fd_sc_hd__and3_1 _6436_ (.A(net188),
    .B(_2408_),
    .C(_2410_),
    .X(_2413_));
 sky130_fd_sc_hd__xnor2_2 _6437_ (.A(_2408_),
    .B(_2412_),
    .Y(_2414_));
 sky130_fd_sc_hd__xnor2_2 _6438_ (.A(_2407_),
    .B(_2414_),
    .Y(_2415_));
 sky130_fd_sc_hd__a31o_1 _6439_ (.A1(net172),
    .A2(_2204_),
    .A3(_2342_),
    .B1(_2341_),
    .X(_2416_));
 sky130_fd_sc_hd__and2_1 _6440_ (.A(_2415_),
    .B(_2416_),
    .X(_2417_));
 sky130_fd_sc_hd__xor2_2 _6441_ (.A(_2415_),
    .B(_2416_),
    .X(_2418_));
 sky130_fd_sc_hd__xnor2_2 _6442_ (.A(_2406_),
    .B(_2418_),
    .Y(_2419_));
 sky130_fd_sc_hd__a21oi_2 _6443_ (.A1(_2332_),
    .A2(_2346_),
    .B1(_2345_),
    .Y(_2420_));
 sky130_fd_sc_hd__or2_1 _6444_ (.A(_2419_),
    .B(_2420_),
    .X(_2421_));
 sky130_fd_sc_hd__xnor2_2 _6445_ (.A(_2419_),
    .B(_2420_),
    .Y(_2422_));
 sky130_fd_sc_hd__xnor2_2 _6446_ (.A(_2399_),
    .B(_2422_),
    .Y(_2423_));
 sky130_fd_sc_hd__a21boi_2 _6447_ (.A1(_2326_),
    .A2(_2350_),
    .B1_N(_2349_),
    .Y(_2424_));
 sky130_fd_sc_hd__nor2_1 _6448_ (.A(_2423_),
    .B(_2424_),
    .Y(_2425_));
 sky130_fd_sc_hd__xor2_2 _6449_ (.A(_2423_),
    .B(_2424_),
    .X(_2426_));
 sky130_fd_sc_hd__xnor2_2 _6450_ (.A(_2389_),
    .B(_2426_),
    .Y(_2427_));
 sky130_fd_sc_hd__a21oi_2 _6451_ (.A1(_2315_),
    .A2(_2354_),
    .B1(_2353_),
    .Y(_2428_));
 sky130_fd_sc_hd__xnor2_2 _6452_ (.A(_2427_),
    .B(_2428_),
    .Y(_2429_));
 sky130_fd_sc_hd__xor2_2 _6453_ (.A(_2314_),
    .B(_2429_),
    .X(_2430_));
 sky130_fd_sc_hd__nor2_1 _6454_ (.A(_2371_),
    .B(_2430_),
    .Y(_2431_));
 sky130_fd_sc_hd__xnor2_2 _6455_ (.A(_2371_),
    .B(_2430_),
    .Y(_2432_));
 sky130_fd_sc_hd__nor2_1 _6456_ (.A(_2361_),
    .B(_2432_),
    .Y(_2433_));
 sky130_fd_sc_hd__xor2_2 _6457_ (.A(_2361_),
    .B(_2432_),
    .X(_2434_));
 sky130_fd_sc_hd__inv_2 _6458_ (.A(_2434_),
    .Y(_2435_));
 sky130_fd_sc_hd__a21o_1 _6459_ (.A1(_2298_),
    .A2(_2365_),
    .B1(_2366_),
    .X(_2436_));
 sky130_fd_sc_hd__a211o_1 _6460_ (.A1(_2290_),
    .A2(_2291_),
    .B1(_2363_),
    .C1(_2289_),
    .X(_2437_));
 sky130_fd_sc_hd__and2_1 _6461_ (.A(_2436_),
    .B(_2437_),
    .X(_2438_));
 sky130_fd_sc_hd__xnor2_1 _6462_ (.A(_2434_),
    .B(_2438_),
    .Y(_2439_));
 sky130_fd_sc_hd__o211ai_1 _6463_ (.A1(_2368_),
    .A2(_2369_),
    .B1(_2294_),
    .C1(_2295_),
    .Y(_2440_));
 sky130_fd_sc_hd__nand2_1 _6464_ (.A(net251),
    .B(_2440_),
    .Y(_2441_));
 sky130_fd_sc_hd__xnor2_1 _6465_ (.A(_2439_),
    .B(_2441_),
    .Y(\mul_la.reg_p[12] ));
 sky130_fd_sc_hd__or2_1 _6466_ (.A(_2439_),
    .B(_2440_),
    .X(_2442_));
 sky130_fd_sc_hd__nand2_1 _6467_ (.A(net251),
    .B(_2442_),
    .Y(_2443_));
 sky130_fd_sc_hd__o21ba_1 _6468_ (.A1(_2435_),
    .A2(_2438_),
    .B1_N(_2433_),
    .X(_2444_));
 sky130_fd_sc_hd__a32oi_4 _6469_ (.A1(_2237_),
    .A2(_2311_),
    .A3(_2388_),
    .B1(_2387_),
    .B2(_2372_),
    .Y(_2445_));
 sky130_fd_sc_hd__a31o_1 _6470_ (.A1(_1756_),
    .A2(_2376_),
    .A3(_2386_),
    .B1(_2385_),
    .X(_2446_));
 sky130_fd_sc_hd__a21bo_1 _6471_ (.A1(_2390_),
    .A2(_2398_),
    .B1_N(_2397_),
    .X(_2447_));
 sky130_fd_sc_hd__a22o_2 _6472_ (.A1(net258),
    .A2(net236),
    .B1(_1610_),
    .B2(net255),
    .X(_2448_));
 sky130_fd_sc_hd__and2_4 _6473_ (.A(_1582_),
    .B(_2448_),
    .X(_2449_));
 sky130_fd_sc_hd__nand2_8 _6474_ (.A(_1582_),
    .B(_2448_),
    .Y(_2450_));
 sky130_fd_sc_hd__or4_2 _6475_ (.A(_1755_),
    .B(_1776_),
    .C(net178),
    .D(_2450_),
    .X(_2451_));
 sky130_fd_sc_hd__a22o_1 _6476_ (.A1(net167),
    .A2(_2376_),
    .B1(_2449_),
    .B2(_1756_),
    .X(_2452_));
 sky130_fd_sc_hd__nand2_1 _6477_ (.A(_2451_),
    .B(_2452_),
    .Y(_2453_));
 sky130_fd_sc_hd__a22o_1 _6478_ (.A1(_1933_),
    .A2(_2175_),
    .B1(_2234_),
    .B2(_1890_),
    .X(_2454_));
 sky130_fd_sc_hd__or4_1 _6479_ (.A(_1891_),
    .B(net169),
    .C(_2176_),
    .D(_2235_),
    .X(_2455_));
 sky130_fd_sc_hd__nor2_1 _6480_ (.A(net170),
    .B(net179),
    .Y(_2456_));
 sky130_fd_sc_hd__and3_1 _6481_ (.A(_2454_),
    .B(_2455_),
    .C(_2456_),
    .X(_2457_));
 sky130_fd_sc_hd__a21oi_1 _6482_ (.A1(_2454_),
    .A2(_2455_),
    .B1(_2456_),
    .Y(_2458_));
 sky130_fd_sc_hd__or2_1 _6483_ (.A(_2457_),
    .B(_2458_),
    .X(_2459_));
 sky130_fd_sc_hd__a31o_1 _6484_ (.A1(net167),
    .A2(_2302_),
    .A3(_2382_),
    .B1(_2381_),
    .X(_2460_));
 sky130_fd_sc_hd__and2b_1 _6485_ (.A_N(_2459_),
    .B(_2460_),
    .X(_2461_));
 sky130_fd_sc_hd__xor2_2 _6486_ (.A(_2459_),
    .B(_2460_),
    .X(_2462_));
 sky130_fd_sc_hd__nor2_1 _6487_ (.A(_2453_),
    .B(_2462_),
    .Y(_2463_));
 sky130_fd_sc_hd__xor2_2 _6488_ (.A(_2453_),
    .B(_2462_),
    .X(_2464_));
 sky130_fd_sc_hd__xnor2_2 _6489_ (.A(_2447_),
    .B(_2464_),
    .Y(_2465_));
 sky130_fd_sc_hd__and2b_1 _6490_ (.A_N(_2465_),
    .B(_2446_),
    .X(_2466_));
 sky130_fd_sc_hd__xnor2_2 _6491_ (.A(_2446_),
    .B(_2465_),
    .Y(_2467_));
 sky130_fd_sc_hd__o31ai_4 _6492_ (.A1(net169),
    .A2(_2115_),
    .A3(_2392_),
    .B1(_2393_),
    .Y(_2468_));
 sky130_fd_sc_hd__o211a_1 _6493_ (.A1(_2022_),
    .A2(_2023_),
    .B1(_2061_),
    .C1(_1700_),
    .X(_2469_));
 sky130_fd_sc_hd__nand2_1 _6494_ (.A(_2005_),
    .B(net183),
    .Y(_2470_));
 sky130_fd_sc_hd__or3_1 _6495_ (.A(_2025_),
    .B(_2062_),
    .C(_2470_),
    .X(_2471_));
 sky130_fd_sc_hd__xor2_1 _6496_ (.A(_2469_),
    .B(_2470_),
    .X(_2472_));
 sky130_fd_sc_hd__nor2_1 _6497_ (.A(net168),
    .B(_2115_),
    .Y(_2473_));
 sky130_fd_sc_hd__xnor2_1 _6498_ (.A(_2472_),
    .B(_2473_),
    .Y(_2474_));
 sky130_fd_sc_hd__o21a_1 _6499_ (.A1(_2402_),
    .A2(_2404_),
    .B1(_2474_),
    .X(_2475_));
 sky130_fd_sc_hd__or3_1 _6500_ (.A(_2402_),
    .B(_2404_),
    .C(_2474_),
    .X(_2476_));
 sky130_fd_sc_hd__and2b_1 _6501_ (.A_N(_2475_),
    .B(_2476_),
    .X(_2477_));
 sky130_fd_sc_hd__xor2_2 _6502_ (.A(_2468_),
    .B(_2477_),
    .X(_2478_));
 sky130_fd_sc_hd__a22o_1 _6503_ (.A1(_1914_),
    .A2(_2204_),
    .B1(_2264_),
    .B2(_1876_),
    .X(_2479_));
 sky130_fd_sc_hd__or4_1 _6504_ (.A(_1877_),
    .B(_1915_),
    .C(_2205_),
    .D(_2265_),
    .X(_2480_));
 sky130_fd_sc_hd__and2_1 _6505_ (.A(_2479_),
    .B(_2480_),
    .X(_2481_));
 sky130_fd_sc_hd__nor2_1 _6506_ (.A(net184),
    .B(net180),
    .Y(_2482_));
 sky130_fd_sc_hd__xor2_2 _6507_ (.A(_2481_),
    .B(_2482_),
    .X(_2483_));
 sky130_fd_sc_hd__nand2_1 _6508_ (.A(net172),
    .B(_2338_),
    .Y(_2484_));
 sky130_fd_sc_hd__a21oi_2 _6509_ (.A1(_1794_),
    .A2(_1802_),
    .B1(_2411_),
    .Y(_2485_));
 sky130_fd_sc_hd__nand2_2 _6510_ (.A(net257),
    .B(net232),
    .Y(_2486_));
 sky130_fd_sc_hd__a21oi_4 _6511_ (.A1(_1732_),
    .A2(_2486_),
    .B1(_1686_),
    .Y(_2487_));
 sky130_fd_sc_hd__a21o_4 _6512_ (.A1(_1732_),
    .A2(_2486_),
    .B1(_1686_),
    .X(_2488_));
 sky130_fd_sc_hd__nand2_1 _6513_ (.A(net187),
    .B(_2487_),
    .Y(_2489_));
 sky130_fd_sc_hd__and3_1 _6514_ (.A(net187),
    .B(_2485_),
    .C(_2487_),
    .X(_2490_));
 sky130_fd_sc_hd__xnor2_2 _6515_ (.A(_2485_),
    .B(_2489_),
    .Y(_2491_));
 sky130_fd_sc_hd__xnor2_2 _6516_ (.A(_2484_),
    .B(_2491_),
    .Y(_2492_));
 sky130_fd_sc_hd__a31o_1 _6517_ (.A1(net172),
    .A2(_2264_),
    .A3(_2414_),
    .B1(_2413_),
    .X(_2493_));
 sky130_fd_sc_hd__and2_1 _6518_ (.A(_2492_),
    .B(_2493_),
    .X(_2494_));
 sky130_fd_sc_hd__xor2_2 _6519_ (.A(_2492_),
    .B(_2493_),
    .X(_2495_));
 sky130_fd_sc_hd__xnor2_2 _6520_ (.A(_2483_),
    .B(_2495_),
    .Y(_2496_));
 sky130_fd_sc_hd__a21o_1 _6521_ (.A1(_2406_),
    .A2(_2418_),
    .B1(_2417_),
    .X(_2497_));
 sky130_fd_sc_hd__nand2b_1 _6522_ (.A_N(_2496_),
    .B(_2497_),
    .Y(_2498_));
 sky130_fd_sc_hd__xnor2_2 _6523_ (.A(_2496_),
    .B(_2497_),
    .Y(_2499_));
 sky130_fd_sc_hd__xor2_2 _6524_ (.A(_2478_),
    .B(_2499_),
    .X(_2500_));
 sky130_fd_sc_hd__o21a_1 _6525_ (.A1(_2399_),
    .A2(_2422_),
    .B1(_2421_),
    .X(_2501_));
 sky130_fd_sc_hd__nand2b_1 _6526_ (.A_N(_2501_),
    .B(_2500_),
    .Y(_2502_));
 sky130_fd_sc_hd__xnor2_2 _6527_ (.A(_2500_),
    .B(_2501_),
    .Y(_2503_));
 sky130_fd_sc_hd__xnor2_2 _6528_ (.A(_2467_),
    .B(_2503_),
    .Y(_2504_));
 sky130_fd_sc_hd__a21oi_2 _6529_ (.A1(_2389_),
    .A2(_2426_),
    .B1(_2425_),
    .Y(_2505_));
 sky130_fd_sc_hd__or2_1 _6530_ (.A(_2504_),
    .B(_2505_),
    .X(_2506_));
 sky130_fd_sc_hd__xor2_2 _6531_ (.A(_2504_),
    .B(_2505_),
    .X(_2507_));
 sky130_fd_sc_hd__nand2b_1 _6532_ (.A_N(_2445_),
    .B(_2507_),
    .Y(_2508_));
 sky130_fd_sc_hd__xnor2_2 _6533_ (.A(_2445_),
    .B(_2507_),
    .Y(_2509_));
 sky130_fd_sc_hd__o32a_1 _6534_ (.A1(_2299_),
    .A2(_2313_),
    .A3(_2429_),
    .B1(_2428_),
    .B2(_2427_),
    .X(_2510_));
 sky130_fd_sc_hd__and2b_1 _6535_ (.A_N(_2510_),
    .B(_2509_),
    .X(_2511_));
 sky130_fd_sc_hd__xnor2_2 _6536_ (.A(_2509_),
    .B(_2510_),
    .Y(_2512_));
 sky130_fd_sc_hd__xor2_2 _6537_ (.A(_2431_),
    .B(_2512_),
    .X(_2513_));
 sky130_fd_sc_hd__xor2_2 _6538_ (.A(_2444_),
    .B(_2513_),
    .X(_2514_));
 sky130_fd_sc_hd__xor2_1 _6539_ (.A(_2443_),
    .B(_2514_),
    .X(\mul_la.reg_p[13] ));
 sky130_fd_sc_hd__a21oi_1 _6540_ (.A1(_2447_),
    .A2(_2464_),
    .B1(_2466_),
    .Y(_2515_));
 sky130_fd_sc_hd__nor2_1 _6541_ (.A(_2451_),
    .B(_2515_),
    .Y(_2516_));
 sky130_fd_sc_hd__xor2_1 _6542_ (.A(_2451_),
    .B(_2515_),
    .X(_2517_));
 sky130_fd_sc_hd__a21o_1 _6543_ (.A1(_2468_),
    .A2(_2476_),
    .B1(_2475_),
    .X(_2518_));
 sky130_fd_sc_hd__a211o_1 _6544_ (.A1(_1766_),
    .A2(_1774_),
    .B1(_2450_),
    .C1(_1725_),
    .X(_2519_));
 sky130_fd_sc_hd__nor2_1 _6545_ (.A(net170),
    .B(net178),
    .Y(_2520_));
 sky130_fd_sc_hd__or3_1 _6546_ (.A(net170),
    .B(net178),
    .C(_2519_),
    .X(_2521_));
 sky130_fd_sc_hd__xnor2_1 _6547_ (.A(_2519_),
    .B(_2520_),
    .Y(_2522_));
 sky130_fd_sc_hd__and2_1 _6548_ (.A(net255),
    .B(net236),
    .X(_2523_));
 sky130_fd_sc_hd__nand2_2 _6549_ (.A(net255),
    .B(net236),
    .Y(_2524_));
 sky130_fd_sc_hd__nor2_1 _6550_ (.A(_1755_),
    .B(net225),
    .Y(_2525_));
 sky130_fd_sc_hd__xnor2_1 _6551_ (.A(_2522_),
    .B(_2525_),
    .Y(_2526_));
 sky130_fd_sc_hd__o211a_2 _6552_ (.A1(_1930_),
    .A2(_1932_),
    .B1(net213),
    .C1(_1720_),
    .X(_2527_));
 sky130_fd_sc_hd__o211a_1 _6553_ (.A1(_1975_),
    .A2(_1977_),
    .B1(net214),
    .C1(_1709_),
    .X(_2528_));
 sky130_fd_sc_hd__or2_1 _6554_ (.A(_2527_),
    .B(_2528_),
    .X(_2529_));
 sky130_fd_sc_hd__and2_1 _6555_ (.A(_2527_),
    .B(_2528_),
    .X(_2530_));
 sky130_fd_sc_hd__xnor2_1 _6556_ (.A(_2527_),
    .B(_2528_),
    .Y(_2531_));
 sky130_fd_sc_hd__nor2_1 _6557_ (.A(_1891_),
    .B(net179),
    .Y(_2532_));
 sky130_fd_sc_hd__xnor2_2 _6558_ (.A(_2531_),
    .B(_2532_),
    .Y(_2533_));
 sky130_fd_sc_hd__a21boi_1 _6559_ (.A1(_2454_),
    .A2(_2456_),
    .B1_N(_2455_),
    .Y(_2534_));
 sky130_fd_sc_hd__nand2b_1 _6560_ (.A_N(_2534_),
    .B(_2533_),
    .Y(_2535_));
 sky130_fd_sc_hd__xnor2_1 _6561_ (.A(_2533_),
    .B(_2534_),
    .Y(_2536_));
 sky130_fd_sc_hd__nand2b_1 _6562_ (.A_N(_2526_),
    .B(_2536_),
    .Y(_2537_));
 sky130_fd_sc_hd__xnor2_1 _6563_ (.A(_2526_),
    .B(_2536_),
    .Y(_2538_));
 sky130_fd_sc_hd__xor2_1 _6564_ (.A(_2518_),
    .B(_2538_),
    .X(_2539_));
 sky130_fd_sc_hd__o21ai_1 _6565_ (.A1(_2461_),
    .A2(_2463_),
    .B1(_2539_),
    .Y(_2540_));
 sky130_fd_sc_hd__or3_1 _6566_ (.A(_2461_),
    .B(_2463_),
    .C(_2539_),
    .X(_2541_));
 sky130_fd_sc_hd__and2_1 _6567_ (.A(_2540_),
    .B(_2541_),
    .X(_2542_));
 sky130_fd_sc_hd__o31a_1 _6568_ (.A1(net168),
    .A2(_2115_),
    .A3(_2472_),
    .B1(_2471_),
    .X(_2543_));
 sky130_fd_sc_hd__a21bo_1 _6569_ (.A1(_2479_),
    .A2(_2482_),
    .B1_N(_2480_),
    .X(_2544_));
 sky130_fd_sc_hd__o2bb2a_1 _6570_ (.A1_N(_2061_),
    .A2_N(net183),
    .B1(net180),
    .B2(_2006_),
    .X(_2545_));
 sky130_fd_sc_hd__and4_1 _6571_ (.A(_2005_),
    .B(_2061_),
    .C(net183),
    .D(_2141_),
    .X(_2546_));
 sky130_fd_sc_hd__or4_1 _6572_ (.A(_2025_),
    .B(_2115_),
    .C(_2545_),
    .D(_2546_),
    .X(_2547_));
 sky130_fd_sc_hd__a2bb2o_1 _6573_ (.A1_N(_2545_),
    .A2_N(_2546_),
    .B1(_2024_),
    .B2(_2116_),
    .X(_2548_));
 sky130_fd_sc_hd__and3_1 _6574_ (.A(_2544_),
    .B(_2547_),
    .C(_2548_),
    .X(_2549_));
 sky130_fd_sc_hd__a21oi_1 _6575_ (.A1(_2547_),
    .A2(_2548_),
    .B1(_2544_),
    .Y(_2550_));
 sky130_fd_sc_hd__or3_1 _6576_ (.A(_2543_),
    .B(_2549_),
    .C(_2550_),
    .X(_2551_));
 sky130_fd_sc_hd__o21ai_1 _6577_ (.A1(_2549_),
    .A2(_2550_),
    .B1(_2543_),
    .Y(_2552_));
 sky130_fd_sc_hd__and2_1 _6578_ (.A(_2551_),
    .B(_2552_),
    .X(_2553_));
 sky130_fd_sc_hd__a22o_1 _6579_ (.A1(_1914_),
    .A2(_2264_),
    .B1(_2338_),
    .B2(_1876_),
    .X(_2554_));
 sky130_fd_sc_hd__or4_1 _6580_ (.A(_1877_),
    .B(_1915_),
    .C(_2265_),
    .D(_2339_),
    .X(_2555_));
 sky130_fd_sc_hd__nor2_1 _6581_ (.A(net184),
    .B(_2205_),
    .Y(_2556_));
 sky130_fd_sc_hd__and3_1 _6582_ (.A(_2554_),
    .B(_2555_),
    .C(_2556_),
    .X(_2557_));
 sky130_fd_sc_hd__a21oi_1 _6583_ (.A1(_2554_),
    .A2(_2555_),
    .B1(_2556_),
    .Y(_2558_));
 sky130_fd_sc_hd__nor2_1 _6584_ (.A(_2557_),
    .B(_2558_),
    .Y(_2559_));
 sky130_fd_sc_hd__nand2_1 _6585_ (.A(net172),
    .B(_2410_),
    .Y(_2560_));
 sky130_fd_sc_hd__a21oi_2 _6586_ (.A1(_1794_),
    .A2(_1802_),
    .B1(_2488_),
    .Y(_2561_));
 sky130_fd_sc_hd__nor2_8 _6587_ (.A(_3372_),
    .B(net233),
    .Y(_2562_));
 sky130_fd_sc_hd__nand2_2 _6588_ (.A(net255),
    .B(_1693_),
    .Y(_2563_));
 sky130_fd_sc_hd__nand2_1 _6589_ (.A(net187),
    .B(_2562_),
    .Y(_2564_));
 sky130_fd_sc_hd__and3_1 _6590_ (.A(net187),
    .B(_2561_),
    .C(_2562_),
    .X(_2565_));
 sky130_fd_sc_hd__xnor2_2 _6591_ (.A(_2561_),
    .B(_2564_),
    .Y(_2566_));
 sky130_fd_sc_hd__xnor2_2 _6592_ (.A(_2560_),
    .B(_2566_),
    .Y(_2567_));
 sky130_fd_sc_hd__a31o_1 _6593_ (.A1(net172),
    .A2(_2338_),
    .A3(_2491_),
    .B1(_2490_),
    .X(_2568_));
 sky130_fd_sc_hd__and2_1 _6594_ (.A(_2567_),
    .B(_2568_),
    .X(_2569_));
 sky130_fd_sc_hd__xor2_2 _6595_ (.A(_2567_),
    .B(_2568_),
    .X(_2570_));
 sky130_fd_sc_hd__xnor2_2 _6596_ (.A(_2559_),
    .B(_2570_),
    .Y(_2571_));
 sky130_fd_sc_hd__a21o_1 _6597_ (.A1(_2483_),
    .A2(_2495_),
    .B1(_2494_),
    .X(_2572_));
 sky130_fd_sc_hd__nand2b_1 _6598_ (.A_N(_2571_),
    .B(_2572_),
    .Y(_2573_));
 sky130_fd_sc_hd__xnor2_2 _6599_ (.A(_2571_),
    .B(_2572_),
    .Y(_2574_));
 sky130_fd_sc_hd__xnor2_2 _6600_ (.A(_2553_),
    .B(_2574_),
    .Y(_2575_));
 sky130_fd_sc_hd__a21bo_1 _6601_ (.A1(_2478_),
    .A2(_2499_),
    .B1_N(_2498_),
    .X(_2576_));
 sky130_fd_sc_hd__and2b_1 _6602_ (.A_N(_2575_),
    .B(_2576_),
    .X(_2577_));
 sky130_fd_sc_hd__xnor2_2 _6603_ (.A(_2575_),
    .B(_2576_),
    .Y(_2578_));
 sky130_fd_sc_hd__xnor2_2 _6604_ (.A(_2542_),
    .B(_2578_),
    .Y(_2579_));
 sky130_fd_sc_hd__a21boi_1 _6605_ (.A1(_2467_),
    .A2(_2503_),
    .B1_N(_2502_),
    .Y(_2580_));
 sky130_fd_sc_hd__nor2_1 _6606_ (.A(_2579_),
    .B(_2580_),
    .Y(_2581_));
 sky130_fd_sc_hd__xor2_1 _6607_ (.A(_2579_),
    .B(_2580_),
    .X(_2582_));
 sky130_fd_sc_hd__xnor2_1 _6608_ (.A(_2517_),
    .B(_2582_),
    .Y(_2583_));
 sky130_fd_sc_hd__a21o_1 _6609_ (.A1(_2506_),
    .A2(_2508_),
    .B1(_2583_),
    .X(_2584_));
 sky130_fd_sc_hd__nand3_1 _6610_ (.A(_2506_),
    .B(_2508_),
    .C(_2583_),
    .Y(_2585_));
 sky130_fd_sc_hd__and2_1 _6611_ (.A(_2584_),
    .B(_2585_),
    .X(_2586_));
 sky130_fd_sc_hd__nand2_1 _6612_ (.A(_2511_),
    .B(_2586_),
    .Y(_2587_));
 sky130_fd_sc_hd__xnor2_2 _6613_ (.A(_2511_),
    .B(_2586_),
    .Y(_2588_));
 sky130_fd_sc_hd__o21ai_1 _6614_ (.A1(_2431_),
    .A2(_2433_),
    .B1(_2512_),
    .Y(_2589_));
 sky130_fd_sc_hd__nand2_1 _6615_ (.A(_2434_),
    .B(_2513_),
    .Y(_2590_));
 sky130_fd_sc_hd__o21a_1 _6616_ (.A1(_2438_),
    .A2(_2590_),
    .B1(_2589_),
    .X(_2591_));
 sky130_fd_sc_hd__xnor2_2 _6617_ (.A(_2588_),
    .B(_2591_),
    .Y(_2592_));
 sky130_fd_sc_hd__and2b_1 _6618_ (.A_N(_2442_),
    .B(_2514_),
    .X(_2593_));
 sky130_fd_sc_hd__nor2_1 _6619_ (.A(_1809_),
    .B(_2593_),
    .Y(_2594_));
 sky130_fd_sc_hd__xnor2_1 _6620_ (.A(_2592_),
    .B(_2594_),
    .Y(\mul_la.reg_p[14] ));
 sky130_fd_sc_hd__a21oi_1 _6621_ (.A1(_2592_),
    .A2(_2593_),
    .B1(_1809_),
    .Y(_2595_));
 sky130_fd_sc_hd__o21ai_1 _6622_ (.A1(_2588_),
    .A2(_2591_),
    .B1(_2587_),
    .Y(_2596_));
 sky130_fd_sc_hd__a21bo_1 _6623_ (.A1(_2518_),
    .A2(_2538_),
    .B1_N(_2540_),
    .X(_2597_));
 sky130_fd_sc_hd__a21bo_1 _6624_ (.A1(_2522_),
    .A2(_2525_),
    .B1_N(_2521_),
    .X(_2598_));
 sky130_fd_sc_hd__and2_1 _6625_ (.A(_2597_),
    .B(_2598_),
    .X(_2599_));
 sky130_fd_sc_hd__inv_2 _6626_ (.A(_2599_),
    .Y(_2600_));
 sky130_fd_sc_hd__xor2_1 _6627_ (.A(_2597_),
    .B(_2598_),
    .X(_2601_));
 sky130_fd_sc_hd__and3_4 _6628_ (.A(net255),
    .B(_1572_),
    .C(_1574_),
    .X(_2602_));
 sky130_fd_sc_hd__nand3_4 _6629_ (.A(net255),
    .B(_1572_),
    .C(_1574_),
    .Y(_2603_));
 sky130_fd_sc_hd__a21o_1 _6630_ (.A1(_1756_),
    .A2(_2602_),
    .B1(_2601_),
    .X(_2604_));
 sky130_fd_sc_hd__nand2_1 _6631_ (.A(_2535_),
    .B(_2537_),
    .Y(_2605_));
 sky130_fd_sc_hd__o21ba_1 _6632_ (.A1(_2543_),
    .A2(_2550_),
    .B1_N(_2549_),
    .X(_2606_));
 sky130_fd_sc_hd__o22a_1 _6633_ (.A1(_1891_),
    .A2(net178),
    .B1(_2450_),
    .B2(net170),
    .X(_2607_));
 sky130_fd_sc_hd__and4b_1 _6634_ (.A_N(net170),
    .B(_1890_),
    .C(_2376_),
    .D(_2449_),
    .X(_2608_));
 sky130_fd_sc_hd__nor2_1 _6635_ (.A(_2607_),
    .B(_2608_),
    .Y(_2609_));
 sky130_fd_sc_hd__nor2_1 _6636_ (.A(_1776_),
    .B(net225),
    .Y(_2610_));
 sky130_fd_sc_hd__xnor2_1 _6637_ (.A(_2609_),
    .B(_2610_),
    .Y(_2611_));
 sky130_fd_sc_hd__o211a_1 _6638_ (.A1(_1975_),
    .A2(_1977_),
    .B1(net213),
    .C1(_1709_),
    .X(_2612_));
 sky130_fd_sc_hd__o211a_1 _6639_ (.A1(_2022_),
    .A2(_2023_),
    .B1(net214),
    .C1(_1700_),
    .X(_2613_));
 sky130_fd_sc_hd__nand2_1 _6640_ (.A(_2612_),
    .B(_2613_),
    .Y(_2614_));
 sky130_fd_sc_hd__xnor2_2 _6641_ (.A(_2612_),
    .B(_2613_),
    .Y(_2615_));
 sky130_fd_sc_hd__nor2_1 _6642_ (.A(net169),
    .B(_2303_),
    .Y(_2616_));
 sky130_fd_sc_hd__xnor2_1 _6643_ (.A(_2615_),
    .B(_2616_),
    .Y(_2617_));
 sky130_fd_sc_hd__a21o_1 _6644_ (.A1(_2529_),
    .A2(_2532_),
    .B1(_2530_),
    .X(_2618_));
 sky130_fd_sc_hd__xor2_1 _6645_ (.A(_2617_),
    .B(_2618_),
    .X(_2619_));
 sky130_fd_sc_hd__and2b_1 _6646_ (.A_N(_2611_),
    .B(_2619_),
    .X(_2620_));
 sky130_fd_sc_hd__xor2_1 _6647_ (.A(_2611_),
    .B(_2619_),
    .X(_2621_));
 sky130_fd_sc_hd__xor2_1 _6648_ (.A(_2606_),
    .B(_2621_),
    .X(_2622_));
 sky130_fd_sc_hd__nand2_1 _6649_ (.A(_2605_),
    .B(_2622_),
    .Y(_2623_));
 sky130_fd_sc_hd__or2_1 _6650_ (.A(_2605_),
    .B(_2622_),
    .X(_2624_));
 sky130_fd_sc_hd__and2_1 _6651_ (.A(_2623_),
    .B(_2624_),
    .X(_2625_));
 sky130_fd_sc_hd__nand2b_1 _6652_ (.A_N(_2546_),
    .B(_2547_),
    .Y(_2626_));
 sky130_fd_sc_hd__a21boi_2 _6653_ (.A1(_2554_),
    .A2(_2556_),
    .B1_N(_2555_),
    .Y(_2627_));
 sky130_fd_sc_hd__a22o_1 _6654_ (.A1(_2061_),
    .A2(_2141_),
    .B1(_2204_),
    .B2(_2005_),
    .X(_2628_));
 sky130_fd_sc_hd__or4_1 _6655_ (.A(_2006_),
    .B(_2062_),
    .C(net180),
    .D(_2205_),
    .X(_2629_));
 sky130_fd_sc_hd__nand2_1 _6656_ (.A(_2628_),
    .B(_2629_),
    .Y(_2630_));
 sky130_fd_sc_hd__and2_1 _6657_ (.A(net182),
    .B(_2116_),
    .X(_2631_));
 sky130_fd_sc_hd__xnor2_2 _6658_ (.A(_2630_),
    .B(_2631_),
    .Y(_2632_));
 sky130_fd_sc_hd__and2b_1 _6659_ (.A_N(_2627_),
    .B(_2632_),
    .X(_2633_));
 sky130_fd_sc_hd__xnor2_2 _6660_ (.A(_2627_),
    .B(_2632_),
    .Y(_2634_));
 sky130_fd_sc_hd__xor2_2 _6661_ (.A(_2626_),
    .B(_2634_),
    .X(_2635_));
 sky130_fd_sc_hd__nand2_1 _6662_ (.A(net186),
    .B(_2338_),
    .Y(_2636_));
 sky130_fd_sc_hd__nor2_1 _6663_ (.A(_1877_),
    .B(_2411_),
    .Y(_2637_));
 sky130_fd_sc_hd__and3_1 _6664_ (.A(net186),
    .B(_2338_),
    .C(_2637_),
    .X(_2638_));
 sky130_fd_sc_hd__xnor2_2 _6665_ (.A(_2636_),
    .B(_2637_),
    .Y(_2639_));
 sky130_fd_sc_hd__nor2_1 _6666_ (.A(net185),
    .B(_2265_),
    .Y(_2640_));
 sky130_fd_sc_hd__xnor2_2 _6667_ (.A(_2639_),
    .B(_2640_),
    .Y(_2641_));
 sky130_fd_sc_hd__nand2_1 _6668_ (.A(net172),
    .B(_2487_),
    .Y(_2642_));
 sky130_fd_sc_hd__and2_4 _6669_ (.A(net255),
    .B(_1694_),
    .X(_2643_));
 sky130_fd_sc_hd__nand2_2 _6670_ (.A(net255),
    .B(_1694_),
    .Y(_2644_));
 sky130_fd_sc_hd__a22o_1 _6671_ (.A1(_1804_),
    .A2(_2562_),
    .B1(_2643_),
    .B2(net187),
    .X(_2645_));
 sky130_fd_sc_hd__nand2b_1 _6672_ (.A_N(_2642_),
    .B(_2645_),
    .Y(_2646_));
 sky130_fd_sc_hd__xor2_2 _6673_ (.A(_2642_),
    .B(_2645_),
    .X(_2647_));
 sky130_fd_sc_hd__a31o_1 _6674_ (.A1(net172),
    .A2(_2410_),
    .A3(_2566_),
    .B1(_2565_),
    .X(_2648_));
 sky130_fd_sc_hd__nand2b_1 _6675_ (.A_N(_2647_),
    .B(_2648_),
    .Y(_2649_));
 sky130_fd_sc_hd__xor2_2 _6676_ (.A(_2647_),
    .B(_2648_),
    .X(_2650_));
 sky130_fd_sc_hd__xnor2_2 _6677_ (.A(_2641_),
    .B(_2650_),
    .Y(_2651_));
 sky130_fd_sc_hd__a21o_1 _6678_ (.A1(_2559_),
    .A2(_2570_),
    .B1(_2569_),
    .X(_2652_));
 sky130_fd_sc_hd__nand2b_1 _6679_ (.A_N(_2651_),
    .B(_2652_),
    .Y(_2653_));
 sky130_fd_sc_hd__xnor2_2 _6680_ (.A(_2651_),
    .B(_2652_),
    .Y(_2654_));
 sky130_fd_sc_hd__xnor2_2 _6681_ (.A(_2635_),
    .B(_2654_),
    .Y(_2655_));
 sky130_fd_sc_hd__a21bo_1 _6682_ (.A1(_2553_),
    .A2(_2574_),
    .B1_N(_2573_),
    .X(_2656_));
 sky130_fd_sc_hd__nand2b_1 _6683_ (.A_N(_2655_),
    .B(_2656_),
    .Y(_2657_));
 sky130_fd_sc_hd__xnor2_2 _6684_ (.A(_2655_),
    .B(_2656_),
    .Y(_2658_));
 sky130_fd_sc_hd__xnor2_2 _6685_ (.A(_2625_),
    .B(_2658_),
    .Y(_2659_));
 sky130_fd_sc_hd__a21oi_2 _6686_ (.A1(_2542_),
    .A2(_2578_),
    .B1(_2577_),
    .Y(_2660_));
 sky130_fd_sc_hd__nor2_1 _6687_ (.A(_2659_),
    .B(_2660_),
    .Y(_2661_));
 sky130_fd_sc_hd__xor2_2 _6688_ (.A(_2659_),
    .B(_2660_),
    .X(_2662_));
 sky130_fd_sc_hd__xnor2_2 _6689_ (.A(_2604_),
    .B(_2662_),
    .Y(_2663_));
 sky130_fd_sc_hd__a21oi_2 _6690_ (.A1(_2517_),
    .A2(_2582_),
    .B1(_2581_),
    .Y(_2664_));
 sky130_fd_sc_hd__nor2_1 _6691_ (.A(_2663_),
    .B(_2664_),
    .Y(_2665_));
 sky130_fd_sc_hd__xor2_2 _6692_ (.A(_2663_),
    .B(_2664_),
    .X(_2666_));
 sky130_fd_sc_hd__xnor2_2 _6693_ (.A(_2516_),
    .B(_2666_),
    .Y(_2667_));
 sky130_fd_sc_hd__xnor2_1 _6694_ (.A(_2584_),
    .B(_2667_),
    .Y(_2668_));
 sky130_fd_sc_hd__xor2_1 _6695_ (.A(_2596_),
    .B(_2668_),
    .X(_2669_));
 sky130_fd_sc_hd__xnor2_1 _6696_ (.A(_2595_),
    .B(_2669_),
    .Y(\mul_la.reg_p[15] ));
 sky130_fd_sc_hd__o21ai_1 _6697_ (.A1(_2606_),
    .A2(_2621_),
    .B1(_2623_),
    .Y(_2670_));
 sky130_fd_sc_hd__a21o_1 _6698_ (.A1(_2609_),
    .A2(_2610_),
    .B1(_2608_),
    .X(_2671_));
 sky130_fd_sc_hd__nand2_1 _6699_ (.A(_2670_),
    .B(_2671_),
    .Y(_2672_));
 sky130_fd_sc_hd__xor2_1 _6700_ (.A(_2670_),
    .B(_2671_),
    .X(_2673_));
 sky130_fd_sc_hd__a21o_1 _6701_ (.A1(net167),
    .A2(_2602_),
    .B1(_2673_),
    .X(_2674_));
 sky130_fd_sc_hd__a21oi_2 _6702_ (.A1(_2617_),
    .A2(_2618_),
    .B1(_2620_),
    .Y(_2675_));
 sky130_fd_sc_hd__a21o_1 _6703_ (.A1(_2626_),
    .A2(_2634_),
    .B1(_2633_),
    .X(_2676_));
 sky130_fd_sc_hd__o22a_1 _6704_ (.A1(_1934_),
    .A2(net178),
    .B1(_2450_),
    .B2(_1891_),
    .X(_2677_));
 sky130_fd_sc_hd__or4_1 _6705_ (.A(_1891_),
    .B(_1934_),
    .C(net178),
    .D(_2450_),
    .X(_2678_));
 sky130_fd_sc_hd__and2b_1 _6706_ (.A_N(_2677_),
    .B(_2678_),
    .X(_2679_));
 sky130_fd_sc_hd__nor2_1 _6707_ (.A(net170),
    .B(net225),
    .Y(_2680_));
 sky130_fd_sc_hd__xnor2_2 _6708_ (.A(_2679_),
    .B(_2680_),
    .Y(_2681_));
 sky130_fd_sc_hd__o211a_1 _6709_ (.A1(_2022_),
    .A2(_2023_),
    .B1(net213),
    .C1(_1700_),
    .X(_2682_));
 sky130_fd_sc_hd__nand2_1 _6710_ (.A(net182),
    .B(net214),
    .Y(_2683_));
 sky130_fd_sc_hd__or3_1 _6711_ (.A(_2025_),
    .B(_2235_),
    .C(_2683_),
    .X(_2684_));
 sky130_fd_sc_hd__xor2_2 _6712_ (.A(_2682_),
    .B(_2683_),
    .X(_2685_));
 sky130_fd_sc_hd__nor2_1 _6713_ (.A(net168),
    .B(net179),
    .Y(_2686_));
 sky130_fd_sc_hd__xnor2_2 _6714_ (.A(_2685_),
    .B(_2686_),
    .Y(_2687_));
 sky130_fd_sc_hd__o31ai_2 _6715_ (.A1(net169),
    .A2(net179),
    .A3(_2615_),
    .B1(_2614_),
    .Y(_2688_));
 sky130_fd_sc_hd__nand2_1 _6716_ (.A(_2687_),
    .B(_2688_),
    .Y(_2689_));
 sky130_fd_sc_hd__nor2_1 _6717_ (.A(_2687_),
    .B(_2688_),
    .Y(_2690_));
 sky130_fd_sc_hd__xor2_1 _6718_ (.A(_2687_),
    .B(_2688_),
    .X(_2691_));
 sky130_fd_sc_hd__xnor2_1 _6719_ (.A(_2681_),
    .B(_2691_),
    .Y(_2692_));
 sky130_fd_sc_hd__nand2_1 _6720_ (.A(_2676_),
    .B(_2692_),
    .Y(_2693_));
 sky130_fd_sc_hd__or2_1 _6721_ (.A(_2676_),
    .B(_2692_),
    .X(_2694_));
 sky130_fd_sc_hd__and2_1 _6722_ (.A(_2693_),
    .B(_2694_),
    .X(_2695_));
 sky130_fd_sc_hd__nand2b_1 _6723_ (.A_N(_2675_),
    .B(_2695_),
    .Y(_2696_));
 sky130_fd_sc_hd__xnor2_2 _6724_ (.A(_2675_),
    .B(_2695_),
    .Y(_2697_));
 sky130_fd_sc_hd__a21bo_1 _6725_ (.A1(_2628_),
    .A2(_2631_),
    .B1_N(_2629_),
    .X(_2698_));
 sky130_fd_sc_hd__a21o_1 _6726_ (.A1(_2639_),
    .A2(_2640_),
    .B1(_2638_),
    .X(_2699_));
 sky130_fd_sc_hd__a22o_1 _6727_ (.A1(_2061_),
    .A2(_2204_),
    .B1(_2264_),
    .B2(_2005_),
    .X(_2700_));
 sky130_fd_sc_hd__or4_1 _6728_ (.A(_2006_),
    .B(_2062_),
    .C(_2205_),
    .D(_2265_),
    .X(_2701_));
 sky130_fd_sc_hd__nand2_1 _6729_ (.A(_2700_),
    .B(_2701_),
    .Y(_2702_));
 sky130_fd_sc_hd__nor2_1 _6730_ (.A(net181),
    .B(net180),
    .Y(_2703_));
 sky130_fd_sc_hd__xnor2_2 _6731_ (.A(_2702_),
    .B(_2703_),
    .Y(_2704_));
 sky130_fd_sc_hd__and2_1 _6732_ (.A(_2699_),
    .B(_2704_),
    .X(_2705_));
 sky130_fd_sc_hd__xor2_2 _6733_ (.A(_2699_),
    .B(_2704_),
    .X(_2706_));
 sky130_fd_sc_hd__xor2_2 _6734_ (.A(_2698_),
    .B(_2706_),
    .X(_2707_));
 sky130_fd_sc_hd__a32oi_2 _6735_ (.A1(_1629_),
    .A2(_1869_),
    .A3(_2487_),
    .B1(_2410_),
    .B2(net186),
    .Y(_2708_));
 sky130_fd_sc_hd__o2111a_1 _6736_ (.A1(_1873_),
    .A2(_1875_),
    .B1(net186),
    .C1(_2410_),
    .D1(_2487_),
    .X(_2709_));
 sky130_fd_sc_hd__nor2_1 _6737_ (.A(_2708_),
    .B(_2709_),
    .Y(_2710_));
 sky130_fd_sc_hd__nand2_1 _6738_ (.A(_1966_),
    .B(_2338_),
    .Y(_2711_));
 sky130_fd_sc_hd__xnor2_2 _6739_ (.A(_2710_),
    .B(_2711_),
    .Y(_2712_));
 sky130_fd_sc_hd__a22o_1 _6740_ (.A1(net172),
    .A2(_2562_),
    .B1(_2643_),
    .B2(_1804_),
    .X(_2713_));
 sky130_fd_sc_hd__nand2_1 _6741_ (.A(_2646_),
    .B(_2713_),
    .Y(_2714_));
 sky130_fd_sc_hd__xnor2_2 _6742_ (.A(_2712_),
    .B(_2714_),
    .Y(_2715_));
 sky130_fd_sc_hd__o21a_1 _6743_ (.A1(_2641_),
    .A2(_2650_),
    .B1(_2649_),
    .X(_2716_));
 sky130_fd_sc_hd__and2b_1 _6744_ (.A_N(_2716_),
    .B(_2715_),
    .X(_2717_));
 sky130_fd_sc_hd__xnor2_2 _6745_ (.A(_2715_),
    .B(_2716_),
    .Y(_2718_));
 sky130_fd_sc_hd__xnor2_2 _6746_ (.A(_2707_),
    .B(_2718_),
    .Y(_2719_));
 sky130_fd_sc_hd__a21bo_1 _6747_ (.A1(_2635_),
    .A2(_2654_),
    .B1_N(_2653_),
    .X(_2720_));
 sky130_fd_sc_hd__nand2b_1 _6748_ (.A_N(_2719_),
    .B(_2720_),
    .Y(_2721_));
 sky130_fd_sc_hd__xnor2_2 _6749_ (.A(_2719_),
    .B(_2720_),
    .Y(_2722_));
 sky130_fd_sc_hd__xnor2_2 _6750_ (.A(_2697_),
    .B(_2722_),
    .Y(_2723_));
 sky130_fd_sc_hd__a21boi_2 _6751_ (.A1(_2625_),
    .A2(_2658_),
    .B1_N(_2657_),
    .Y(_2724_));
 sky130_fd_sc_hd__nor2_1 _6752_ (.A(_2723_),
    .B(_2724_),
    .Y(_2725_));
 sky130_fd_sc_hd__xor2_2 _6753_ (.A(_2723_),
    .B(_2724_),
    .X(_2726_));
 sky130_fd_sc_hd__xnor2_2 _6754_ (.A(_2674_),
    .B(_2726_),
    .Y(_2727_));
 sky130_fd_sc_hd__a21oi_2 _6755_ (.A1(_2604_),
    .A2(_2662_),
    .B1(_2661_),
    .Y(_2728_));
 sky130_fd_sc_hd__or2_1 _6756_ (.A(_2727_),
    .B(_2728_),
    .X(_2729_));
 sky130_fd_sc_hd__xnor2_2 _6757_ (.A(_2727_),
    .B(_2728_),
    .Y(_2730_));
 sky130_fd_sc_hd__xnor2_2 _6758_ (.A(_2600_),
    .B(_2730_),
    .Y(_2731_));
 sky130_fd_sc_hd__a21oi_2 _6759_ (.A1(_2516_),
    .A2(_2666_),
    .B1(_2665_),
    .Y(_2732_));
 sky130_fd_sc_hd__or2_1 _6760_ (.A(_2731_),
    .B(_2732_),
    .X(_2733_));
 sky130_fd_sc_hd__nand2_1 _6761_ (.A(_2731_),
    .B(_2732_),
    .Y(_2734_));
 sky130_fd_sc_hd__and2_1 _6762_ (.A(_2733_),
    .B(_2734_),
    .X(_2735_));
 sky130_fd_sc_hd__xnor2_1 _6763_ (.A(_2731_),
    .B(_2732_),
    .Y(_2736_));
 sky130_fd_sc_hd__a21o_1 _6764_ (.A1(_2584_),
    .A2(_2587_),
    .B1(_2667_),
    .X(_2737_));
 sky130_fd_sc_hd__or3_2 _6765_ (.A(_2588_),
    .B(_2589_),
    .C(_2668_),
    .X(_2738_));
 sky130_fd_sc_hd__a2111o_2 _6766_ (.A1(_2436_),
    .A2(_2437_),
    .B1(_2588_),
    .C1(_2590_),
    .D1(_2668_),
    .X(_2739_));
 sky130_fd_sc_hd__nand3_4 _6767_ (.A(_2737_),
    .B(_2738_),
    .C(_2739_),
    .Y(_2740_));
 sky130_fd_sc_hd__xnor2_2 _6768_ (.A(_2735_),
    .B(_2740_),
    .Y(_2741_));
 sky130_fd_sc_hd__and3_1 _6769_ (.A(_2592_),
    .B(_2593_),
    .C(_2669_),
    .X(_2742_));
 sky130_fd_sc_hd__nor2_1 _6770_ (.A(_1809_),
    .B(_2742_),
    .Y(_2743_));
 sky130_fd_sc_hd__xnor2_1 _6771_ (.A(_2741_),
    .B(_2743_),
    .Y(\mul_la.reg_p[16] ));
 sky130_fd_sc_hd__o21ai_2 _6772_ (.A1(_2600_),
    .A2(_2730_),
    .B1(_2729_),
    .Y(_2744_));
 sky130_fd_sc_hd__o31a_1 _6773_ (.A1(net170),
    .A2(_2524_),
    .A3(_2677_),
    .B1(_2678_),
    .X(_2745_));
 sky130_fd_sc_hd__a21oi_2 _6774_ (.A1(_2693_),
    .A2(_2696_),
    .B1(_2745_),
    .Y(_2746_));
 sky130_fd_sc_hd__a21o_1 _6775_ (.A1(_2693_),
    .A2(_2696_),
    .B1(_2745_),
    .X(_2747_));
 sky130_fd_sc_hd__and3_1 _6776_ (.A(_2693_),
    .B(_2696_),
    .C(_2745_),
    .X(_2748_));
 sky130_fd_sc_hd__o22ai_4 _6777_ (.A1(net170),
    .A2(_2603_),
    .B1(_2746_),
    .B2(_2748_),
    .Y(_2749_));
 sky130_fd_sc_hd__o21ai_2 _6778_ (.A1(_2681_),
    .A2(_2690_),
    .B1(_2689_),
    .Y(_2750_));
 sky130_fd_sc_hd__a21o_1 _6779_ (.A1(_2698_),
    .A2(_2706_),
    .B1(_2705_),
    .X(_2751_));
 sky130_fd_sc_hd__a22o_1 _6780_ (.A1(_1978_),
    .A2(_2376_),
    .B1(_2449_),
    .B2(_1933_),
    .X(_2752_));
 sky130_fd_sc_hd__or4_1 _6781_ (.A(net169),
    .B(net168),
    .C(net178),
    .D(_2450_),
    .X(_2753_));
 sky130_fd_sc_hd__nand2_1 _6782_ (.A(_2752_),
    .B(_2753_),
    .Y(_2754_));
 sky130_fd_sc_hd__nor2_1 _6783_ (.A(_1891_),
    .B(net225),
    .Y(_2755_));
 sky130_fd_sc_hd__xnor2_2 _6784_ (.A(_2754_),
    .B(_2755_),
    .Y(_2756_));
 sky130_fd_sc_hd__a22o_1 _6785_ (.A1(_2141_),
    .A2(net214),
    .B1(net213),
    .B2(net182),
    .X(_2757_));
 sky130_fd_sc_hd__and4_1 _6786_ (.A(net182),
    .B(_2141_),
    .C(net214),
    .D(net213),
    .X(_2758_));
 sky130_fd_sc_hd__nand4_1 _6787_ (.A(net182),
    .B(_2141_),
    .C(net214),
    .D(net213),
    .Y(_2759_));
 sky130_fd_sc_hd__or4b_1 _6788_ (.A(_2025_),
    .B(_2758_),
    .C(net179),
    .D_N(_2757_),
    .X(_2760_));
 sky130_fd_sc_hd__a22o_1 _6789_ (.A1(_2024_),
    .A2(_2302_),
    .B1(_2757_),
    .B2(_2759_),
    .X(_2761_));
 sky130_fd_sc_hd__nand2_1 _6790_ (.A(_2760_),
    .B(_2761_),
    .Y(_2762_));
 sky130_fd_sc_hd__o31a_1 _6791_ (.A1(net168),
    .A2(net179),
    .A3(_2685_),
    .B1(_2684_),
    .X(_2763_));
 sky130_fd_sc_hd__nor2_1 _6792_ (.A(_2762_),
    .B(_2763_),
    .Y(_2764_));
 sky130_fd_sc_hd__nand2_1 _6793_ (.A(_2762_),
    .B(_2763_),
    .Y(_2765_));
 sky130_fd_sc_hd__and2b_1 _6794_ (.A_N(_2764_),
    .B(_2765_),
    .X(_2766_));
 sky130_fd_sc_hd__xnor2_2 _6795_ (.A(_2756_),
    .B(_2766_),
    .Y(_2767_));
 sky130_fd_sc_hd__and2b_1 _6796_ (.A_N(_2767_),
    .B(_2751_),
    .X(_2768_));
 sky130_fd_sc_hd__xnor2_2 _6797_ (.A(_2751_),
    .B(_2767_),
    .Y(_2769_));
 sky130_fd_sc_hd__xnor2_2 _6798_ (.A(_2750_),
    .B(_2769_),
    .Y(_2770_));
 sky130_fd_sc_hd__a21bo_1 _6799_ (.A1(_2700_),
    .A2(_2703_),
    .B1_N(_2701_),
    .X(_2771_));
 sky130_fd_sc_hd__o21bai_1 _6800_ (.A1(_2708_),
    .A2(_2711_),
    .B1_N(_2709_),
    .Y(_2772_));
 sky130_fd_sc_hd__a22o_1 _6801_ (.A1(_2061_),
    .A2(_2264_),
    .B1(_2338_),
    .B2(_2005_),
    .X(_2773_));
 sky130_fd_sc_hd__or4_1 _6802_ (.A(_2006_),
    .B(_2062_),
    .C(_2265_),
    .D(_2339_),
    .X(_2774_));
 sky130_fd_sc_hd__nor2_1 _6803_ (.A(net181),
    .B(_2205_),
    .Y(_2775_));
 sky130_fd_sc_hd__nand3_1 _6804_ (.A(_2773_),
    .B(_2774_),
    .C(_2775_),
    .Y(_2776_));
 sky130_fd_sc_hd__a21o_1 _6805_ (.A1(_2773_),
    .A2(_2774_),
    .B1(_2775_),
    .X(_2777_));
 sky130_fd_sc_hd__nand3_1 _6806_ (.A(_2772_),
    .B(_2776_),
    .C(_2777_),
    .Y(_2778_));
 sky130_fd_sc_hd__a21o_1 _6807_ (.A1(_2776_),
    .A2(_2777_),
    .B1(_2772_),
    .X(_2779_));
 sky130_fd_sc_hd__and3_1 _6808_ (.A(_2771_),
    .B(_2778_),
    .C(_2779_),
    .X(_2780_));
 sky130_fd_sc_hd__a21oi_1 _6809_ (.A1(_2778_),
    .A2(_2779_),
    .B1(_2771_),
    .Y(_2781_));
 sky130_fd_sc_hd__a32o_1 _6810_ (.A1(_1629_),
    .A2(_1869_),
    .A3(_2562_),
    .B1(_2487_),
    .B2(net186),
    .X(_2782_));
 sky130_fd_sc_hd__o2111a_1 _6811_ (.A1(_1873_),
    .A2(_1875_),
    .B1(net186),
    .C1(_2487_),
    .D1(_2562_),
    .X(_2783_));
 sky130_fd_sc_hd__or4_1 _6812_ (.A(_1877_),
    .B(_1915_),
    .C(_2488_),
    .D(_2563_),
    .X(_2784_));
 sky130_fd_sc_hd__nor2_1 _6813_ (.A(net185),
    .B(_2411_),
    .Y(_2785_));
 sky130_fd_sc_hd__a21oi_1 _6814_ (.A1(_2782_),
    .A2(_2784_),
    .B1(_2785_),
    .Y(_2786_));
 sky130_fd_sc_hd__and3_1 _6815_ (.A(_2782_),
    .B(_2784_),
    .C(_2785_),
    .X(_2787_));
 sky130_fd_sc_hd__a2bb2o_1 _6816_ (.A1_N(_2786_),
    .A2_N(_2787_),
    .B1(net172),
    .B2(_2643_),
    .X(_2788_));
 sky130_fd_sc_hd__a21bo_1 _6817_ (.A1(_2712_),
    .A2(_2713_),
    .B1_N(_2646_),
    .X(_2789_));
 sky130_fd_sc_hd__nand2_1 _6818_ (.A(_2788_),
    .B(_2789_),
    .Y(_2790_));
 sky130_fd_sc_hd__xnor2_1 _6819_ (.A(_2788_),
    .B(_2789_),
    .Y(_2791_));
 sky130_fd_sc_hd__or3_2 _6820_ (.A(_2780_),
    .B(_2781_),
    .C(_2791_),
    .X(_2792_));
 sky130_fd_sc_hd__o21ai_1 _6821_ (.A1(_2780_),
    .A2(_2781_),
    .B1(_2791_),
    .Y(_2793_));
 sky130_fd_sc_hd__nand2_2 _6822_ (.A(_2792_),
    .B(_2793_),
    .Y(_2794_));
 sky130_fd_sc_hd__a21oi_2 _6823_ (.A1(_2707_),
    .A2(_2718_),
    .B1(_2717_),
    .Y(_2795_));
 sky130_fd_sc_hd__or2_1 _6824_ (.A(_2794_),
    .B(_2795_),
    .X(_2796_));
 sky130_fd_sc_hd__xnor2_2 _6825_ (.A(_2794_),
    .B(_2795_),
    .Y(_2797_));
 sky130_fd_sc_hd__xnor2_2 _6826_ (.A(_2770_),
    .B(_2797_),
    .Y(_2798_));
 sky130_fd_sc_hd__a21boi_2 _6827_ (.A1(_2697_),
    .A2(_2722_),
    .B1_N(_2721_),
    .Y(_2799_));
 sky130_fd_sc_hd__nor2_1 _6828_ (.A(_2798_),
    .B(_2799_),
    .Y(_2800_));
 sky130_fd_sc_hd__xor2_2 _6829_ (.A(_2798_),
    .B(_2799_),
    .X(_2801_));
 sky130_fd_sc_hd__xnor2_2 _6830_ (.A(_2749_),
    .B(_2801_),
    .Y(_2802_));
 sky130_fd_sc_hd__a21oi_2 _6831_ (.A1(_2674_),
    .A2(_2726_),
    .B1(_2725_),
    .Y(_2803_));
 sky130_fd_sc_hd__or2_1 _6832_ (.A(_2802_),
    .B(_2803_),
    .X(_2804_));
 sky130_fd_sc_hd__xnor2_2 _6833_ (.A(_2802_),
    .B(_2803_),
    .Y(_2805_));
 sky130_fd_sc_hd__xor2_2 _6834_ (.A(_2672_),
    .B(_2805_),
    .X(_2806_));
 sky130_fd_sc_hd__and2_1 _6835_ (.A(_2744_),
    .B(_2806_),
    .X(_2807_));
 sky130_fd_sc_hd__nand2_1 _6836_ (.A(_2744_),
    .B(_2806_),
    .Y(_2808_));
 sky130_fd_sc_hd__nor2_1 _6837_ (.A(_2744_),
    .B(_2806_),
    .Y(_2809_));
 sky130_fd_sc_hd__nor2_1 _6838_ (.A(_2807_),
    .B(_2809_),
    .Y(_2810_));
 sky130_fd_sc_hd__xnor2_1 _6839_ (.A(_2744_),
    .B(_2806_),
    .Y(_2811_));
 sky130_fd_sc_hd__a21bo_1 _6840_ (.A1(_2735_),
    .A2(_2740_),
    .B1_N(_2733_),
    .X(_2812_));
 sky130_fd_sc_hd__xnor2_2 _6841_ (.A(_2810_),
    .B(_2812_),
    .Y(_2813_));
 sky130_fd_sc_hd__a21o_1 _6842_ (.A1(_2741_),
    .A2(_2742_),
    .B1(_1809_),
    .X(_2814_));
 sky130_fd_sc_hd__xor2_1 _6843_ (.A(_2813_),
    .B(_2814_),
    .X(\mul_la.reg_p[17] ));
 sky130_fd_sc_hd__a21o_1 _6844_ (.A1(_2750_),
    .A2(_2769_),
    .B1(_2768_),
    .X(_2815_));
 sky130_fd_sc_hd__a21bo_1 _6845_ (.A1(_2752_),
    .A2(_2755_),
    .B1_N(_2753_),
    .X(_2816_));
 sky130_fd_sc_hd__nand2_1 _6846_ (.A(_2815_),
    .B(_2816_),
    .Y(_2817_));
 sky130_fd_sc_hd__or2_1 _6847_ (.A(_2815_),
    .B(_2816_),
    .X(_2818_));
 sky130_fd_sc_hd__a22o_1 _6848_ (.A1(_1890_),
    .A2(_2602_),
    .B1(_2817_),
    .B2(_2818_),
    .X(_2819_));
 sky130_fd_sc_hd__a21o_1 _6849_ (.A1(_2756_),
    .A2(_2766_),
    .B1(_2764_),
    .X(_2820_));
 sky130_fd_sc_hd__a21boi_1 _6850_ (.A1(_2771_),
    .A2(_2779_),
    .B1_N(_2778_),
    .Y(_2821_));
 sky130_fd_sc_hd__o211a_1 _6851_ (.A1(_1975_),
    .A2(_1977_),
    .B1(_2449_),
    .C1(_1709_),
    .X(_2822_));
 sky130_fd_sc_hd__o211a_1 _6852_ (.A1(_2022_),
    .A2(_2023_),
    .B1(_2376_),
    .C1(_1700_),
    .X(_2823_));
 sky130_fd_sc_hd__nand2_1 _6853_ (.A(_2822_),
    .B(_2823_),
    .Y(_2824_));
 sky130_fd_sc_hd__xnor2_1 _6854_ (.A(_2822_),
    .B(_2823_),
    .Y(_2825_));
 sky130_fd_sc_hd__nor2_1 _6855_ (.A(net169),
    .B(net225),
    .Y(_2826_));
 sky130_fd_sc_hd__xnor2_1 _6856_ (.A(_2825_),
    .B(_2826_),
    .Y(_2827_));
 sky130_fd_sc_hd__o311a_1 _6857_ (.A1(_2133_),
    .A2(_2134_),
    .A3(_2140_),
    .B1(net213),
    .C1(_1672_),
    .X(_2828_));
 sky130_fd_sc_hd__o211a_1 _6858_ (.A1(_2201_),
    .A2(_2203_),
    .B1(_1670_),
    .C1(net214),
    .X(_2829_));
 sky130_fd_sc_hd__and2_1 _6859_ (.A(_2828_),
    .B(_2829_),
    .X(_2830_));
 sky130_fd_sc_hd__xnor2_1 _6860_ (.A(_2828_),
    .B(_2829_),
    .Y(_2831_));
 sky130_fd_sc_hd__nand2_1 _6861_ (.A(net182),
    .B(_2302_),
    .Y(_2832_));
 sky130_fd_sc_hd__xor2_1 _6862_ (.A(_2831_),
    .B(_2832_),
    .X(_2833_));
 sky130_fd_sc_hd__a31o_1 _6863_ (.A1(_2024_),
    .A2(_2302_),
    .A3(_2757_),
    .B1(_2758_),
    .X(_2834_));
 sky130_fd_sc_hd__and2_1 _6864_ (.A(_2833_),
    .B(_2834_),
    .X(_2835_));
 sky130_fd_sc_hd__xor2_1 _6865_ (.A(_2833_),
    .B(_2834_),
    .X(_2836_));
 sky130_fd_sc_hd__xnor2_1 _6866_ (.A(_2827_),
    .B(_2836_),
    .Y(_2837_));
 sky130_fd_sc_hd__nor2_1 _6867_ (.A(_2821_),
    .B(_2837_),
    .Y(_2838_));
 sky130_fd_sc_hd__and2_1 _6868_ (.A(_2821_),
    .B(_2837_),
    .X(_2839_));
 sky130_fd_sc_hd__or2_1 _6869_ (.A(_2838_),
    .B(_2839_),
    .X(_2840_));
 sky130_fd_sc_hd__and2b_1 _6870_ (.A_N(_2840_),
    .B(_2820_),
    .X(_2841_));
 sky130_fd_sc_hd__xnor2_1 _6871_ (.A(_2820_),
    .B(_2840_),
    .Y(_2842_));
 sky130_fd_sc_hd__a32o_1 _6872_ (.A1(_1629_),
    .A2(_1869_),
    .A3(_2643_),
    .B1(_2562_),
    .B2(net186),
    .X(_2843_));
 sky130_fd_sc_hd__or3b_1 _6873_ (.A(net185),
    .B(_2488_),
    .C_N(_2843_),
    .X(_2844_));
 sky130_fd_sc_hd__a21o_1 _6874_ (.A1(_1966_),
    .A2(_2487_),
    .B1(_2843_),
    .X(_2845_));
 sky130_fd_sc_hd__and2_1 _6875_ (.A(_2844_),
    .B(_2845_),
    .X(_2846_));
 sky130_fd_sc_hd__nand2_1 _6876_ (.A(_2774_),
    .B(_2776_),
    .Y(_2847_));
 sky130_fd_sc_hd__a21o_1 _6877_ (.A1(_2782_),
    .A2(_2785_),
    .B1(_2783_),
    .X(_2848_));
 sky130_fd_sc_hd__a22o_1 _6878_ (.A1(_2061_),
    .A2(_2338_),
    .B1(_2410_),
    .B2(_2005_),
    .X(_2849_));
 sky130_fd_sc_hd__or4_1 _6879_ (.A(_2006_),
    .B(_2062_),
    .C(_2339_),
    .D(_2411_),
    .X(_2850_));
 sky130_fd_sc_hd__nor2_1 _6880_ (.A(net181),
    .B(_2265_),
    .Y(_2851_));
 sky130_fd_sc_hd__nand3_1 _6881_ (.A(_2849_),
    .B(_2850_),
    .C(_2851_),
    .Y(_2852_));
 sky130_fd_sc_hd__a21o_1 _6882_ (.A1(_2849_),
    .A2(_2850_),
    .B1(_2851_),
    .X(_2853_));
 sky130_fd_sc_hd__nand3_1 _6883_ (.A(_2848_),
    .B(_2852_),
    .C(_2853_),
    .Y(_2854_));
 sky130_fd_sc_hd__a21o_1 _6884_ (.A1(_2852_),
    .A2(_2853_),
    .B1(_2848_),
    .X(_2855_));
 sky130_fd_sc_hd__and3_1 _6885_ (.A(_2847_),
    .B(_2854_),
    .C(_2855_),
    .X(_2856_));
 sky130_fd_sc_hd__a21oi_1 _6886_ (.A1(_2854_),
    .A2(_2855_),
    .B1(_2847_),
    .Y(_2857_));
 sky130_fd_sc_hd__nor3b_2 _6887_ (.A(_2856_),
    .B(_2857_),
    .C_N(_2846_),
    .Y(_2858_));
 sky130_fd_sc_hd__o21ba_1 _6888_ (.A1(_2856_),
    .A2(_2857_),
    .B1_N(_2846_),
    .X(_2859_));
 sky130_fd_sc_hd__a211o_1 _6889_ (.A1(_2790_),
    .A2(_2792_),
    .B1(_2858_),
    .C1(_2859_),
    .X(_2860_));
 sky130_fd_sc_hd__o211ai_2 _6890_ (.A1(_2858_),
    .A2(_2859_),
    .B1(_2790_),
    .C1(_2792_),
    .Y(_2861_));
 sky130_fd_sc_hd__and3_1 _6891_ (.A(_2842_),
    .B(_2860_),
    .C(_2861_),
    .X(_2862_));
 sky130_fd_sc_hd__a21oi_1 _6892_ (.A1(_2860_),
    .A2(_2861_),
    .B1(_2842_),
    .Y(_2863_));
 sky130_fd_sc_hd__nor2_1 _6893_ (.A(_2862_),
    .B(_2863_),
    .Y(_2864_));
 sky130_fd_sc_hd__o21ai_2 _6894_ (.A1(_2770_),
    .A2(_2797_),
    .B1(_2796_),
    .Y(_2865_));
 sky130_fd_sc_hd__and2_1 _6895_ (.A(_2864_),
    .B(_2865_),
    .X(_2866_));
 sky130_fd_sc_hd__xor2_2 _6896_ (.A(_2864_),
    .B(_2865_),
    .X(_2867_));
 sky130_fd_sc_hd__xnor2_2 _6897_ (.A(_2819_),
    .B(_2867_),
    .Y(_2868_));
 sky130_fd_sc_hd__a21oi_2 _6898_ (.A1(_2749_),
    .A2(_2801_),
    .B1(_2800_),
    .Y(_2869_));
 sky130_fd_sc_hd__or2_1 _6899_ (.A(_2868_),
    .B(_2869_),
    .X(_2870_));
 sky130_fd_sc_hd__xnor2_2 _6900_ (.A(_2868_),
    .B(_2869_),
    .Y(_2871_));
 sky130_fd_sc_hd__xnor2_2 _6901_ (.A(_2746_),
    .B(_2871_),
    .Y(_2872_));
 sky130_fd_sc_hd__o21a_1 _6902_ (.A1(_2672_),
    .A2(_2805_),
    .B1(_2804_),
    .X(_2873_));
 sky130_fd_sc_hd__and2b_1 _6903_ (.A_N(_2873_),
    .B(_2872_),
    .X(_2874_));
 sky130_fd_sc_hd__xor2_2 _6904_ (.A(_2872_),
    .B(_2873_),
    .X(_2875_));
 sky130_fd_sc_hd__inv_2 _6905_ (.A(_2875_),
    .Y(_2876_));
 sky130_fd_sc_hd__a21oi_1 _6906_ (.A1(_2733_),
    .A2(_2808_),
    .B1(_2809_),
    .Y(_2877_));
 sky130_fd_sc_hd__a31o_1 _6907_ (.A1(_2735_),
    .A2(_2740_),
    .A3(_2810_),
    .B1(_2877_),
    .X(_2878_));
 sky130_fd_sc_hd__xnor2_2 _6908_ (.A(_2876_),
    .B(_2878_),
    .Y(_2879_));
 sky130_fd_sc_hd__and2_1 _6909_ (.A(_2741_),
    .B(_2813_),
    .X(_2880_));
 sky130_fd_sc_hd__a21oi_1 _6910_ (.A1(_2742_),
    .A2(_2880_),
    .B1(_1809_),
    .Y(_2881_));
 sky130_fd_sc_hd__xnor2_1 _6911_ (.A(_2879_),
    .B(_2881_),
    .Y(\mul_la.reg_p[18] ));
 sky130_fd_sc_hd__a31o_1 _6912_ (.A1(_2742_),
    .A2(_2879_),
    .A3(_2880_),
    .B1(_1809_),
    .X(_2882_));
 sky130_fd_sc_hd__o21ai_4 _6913_ (.A1(_2747_),
    .A2(_2871_),
    .B1(_2870_),
    .Y(_2883_));
 sky130_fd_sc_hd__o31a_1 _6914_ (.A1(net169),
    .A2(net225),
    .A3(_2825_),
    .B1(_2824_),
    .X(_2884_));
 sky130_fd_sc_hd__o21bai_2 _6915_ (.A1(_2838_),
    .A2(_2841_),
    .B1_N(_2884_),
    .Y(_2885_));
 sky130_fd_sc_hd__or3b_1 _6916_ (.A(_2838_),
    .B(_2841_),
    .C_N(_2884_),
    .X(_2886_));
 sky130_fd_sc_hd__o2bb2a_1 _6917_ (.A1_N(_2885_),
    .A2_N(_2886_),
    .B1(net169),
    .B2(_2603_),
    .X(_2887_));
 sky130_fd_sc_hd__a22o_1 _6918_ (.A1(_1966_),
    .A2(_2562_),
    .B1(_2643_),
    .B2(net186),
    .X(_2888_));
 sky130_fd_sc_hd__nand2_1 _6919_ (.A(_2850_),
    .B(_2852_),
    .Y(_2889_));
 sky130_fd_sc_hd__a211o_1 _6920_ (.A1(_2055_),
    .A2(net215),
    .B1(_2411_),
    .C1(_1618_),
    .X(_2890_));
 sky130_fd_sc_hd__o211a_1 _6921_ (.A1(_2003_),
    .A2(_2004_),
    .B1(_2487_),
    .C1(_1621_),
    .X(_2891_));
 sky130_fd_sc_hd__xor2_1 _6922_ (.A(_2890_),
    .B(_2891_),
    .X(_2892_));
 sky130_fd_sc_hd__or2_1 _6923_ (.A(net181),
    .B(_2339_),
    .X(_2893_));
 sky130_fd_sc_hd__nor2_1 _6924_ (.A(_2892_),
    .B(_2893_),
    .Y(_2894_));
 sky130_fd_sc_hd__xnor2_1 _6925_ (.A(_2892_),
    .B(_2893_),
    .Y(_2895_));
 sky130_fd_sc_hd__nor2_1 _6926_ (.A(_2844_),
    .B(_2895_),
    .Y(_2896_));
 sky130_fd_sc_hd__xor2_1 _6927_ (.A(_2844_),
    .B(_2895_),
    .X(_2897_));
 sky130_fd_sc_hd__xor2_1 _6928_ (.A(_2889_),
    .B(_2897_),
    .X(_2898_));
 sky130_fd_sc_hd__and2_1 _6929_ (.A(_2888_),
    .B(_2898_),
    .X(_2899_));
 sky130_fd_sc_hd__xor2_1 _6930_ (.A(_2888_),
    .B(_2898_),
    .X(_2900_));
 sky130_fd_sc_hd__nand2_1 _6931_ (.A(_2858_),
    .B(_2900_),
    .Y(_2901_));
 sky130_fd_sc_hd__xnor2_1 _6932_ (.A(_2858_),
    .B(_2900_),
    .Y(_2902_));
 sky130_fd_sc_hd__a21o_1 _6933_ (.A1(_2827_),
    .A2(_2836_),
    .B1(_2835_),
    .X(_2903_));
 sky130_fd_sc_hd__a21boi_1 _6934_ (.A1(_2847_),
    .A2(_2855_),
    .B1_N(_2854_),
    .Y(_2904_));
 sky130_fd_sc_hd__o211a_1 _6935_ (.A1(_2022_),
    .A2(_2023_),
    .B1(_2449_),
    .C1(_1700_),
    .X(_2905_));
 sky130_fd_sc_hd__nand2_1 _6936_ (.A(net182),
    .B(_2376_),
    .Y(_2906_));
 sky130_fd_sc_hd__or3_1 _6937_ (.A(_2025_),
    .B(_2450_),
    .C(_2906_),
    .X(_2907_));
 sky130_fd_sc_hd__xor2_2 _6938_ (.A(_2905_),
    .B(_2906_),
    .X(_2908_));
 sky130_fd_sc_hd__nor2_1 _6939_ (.A(net168),
    .B(net225),
    .Y(_2909_));
 sky130_fd_sc_hd__xnor2_2 _6940_ (.A(_2908_),
    .B(_2909_),
    .Y(_2910_));
 sky130_fd_sc_hd__o211a_1 _6941_ (.A1(_2201_),
    .A2(_2203_),
    .B1(net213),
    .C1(_1670_),
    .X(_2911_));
 sky130_fd_sc_hd__o211a_1 _6942_ (.A1(_2260_),
    .A2(_2263_),
    .B1(_1676_),
    .C1(net214),
    .X(_2912_));
 sky130_fd_sc_hd__nand2_1 _6943_ (.A(_2911_),
    .B(_2912_),
    .Y(_2913_));
 sky130_fd_sc_hd__xnor2_2 _6944_ (.A(_2911_),
    .B(_2912_),
    .Y(_2914_));
 sky130_fd_sc_hd__nor2_1 _6945_ (.A(_2142_),
    .B(net179),
    .Y(_2915_));
 sky130_fd_sc_hd__xnor2_1 _6946_ (.A(_2914_),
    .B(_2915_),
    .Y(_2916_));
 sky130_fd_sc_hd__o21bai_1 _6947_ (.A1(_2831_),
    .A2(_2832_),
    .B1_N(_2830_),
    .Y(_2917_));
 sky130_fd_sc_hd__and2_1 _6948_ (.A(_2916_),
    .B(_2917_),
    .X(_2918_));
 sky130_fd_sc_hd__xor2_1 _6949_ (.A(_2916_),
    .B(_2917_),
    .X(_2919_));
 sky130_fd_sc_hd__xor2_1 _6950_ (.A(_2910_),
    .B(_2919_),
    .X(_2920_));
 sky130_fd_sc_hd__and2b_1 _6951_ (.A_N(_2904_),
    .B(_2920_),
    .X(_2921_));
 sky130_fd_sc_hd__xnor2_1 _6952_ (.A(_2904_),
    .B(_2920_),
    .Y(_2922_));
 sky130_fd_sc_hd__and2_1 _6953_ (.A(_2903_),
    .B(_2922_),
    .X(_2923_));
 sky130_fd_sc_hd__xor2_1 _6954_ (.A(_2903_),
    .B(_2922_),
    .X(_2924_));
 sky130_fd_sc_hd__nand2b_1 _6955_ (.A_N(_2902_),
    .B(_2924_),
    .Y(_2925_));
 sky130_fd_sc_hd__xnor2_1 _6956_ (.A(_2902_),
    .B(_2924_),
    .Y(_2926_));
 sky130_fd_sc_hd__a21bo_1 _6957_ (.A1(_2842_),
    .A2(_2861_),
    .B1_N(_2860_),
    .X(_2927_));
 sky130_fd_sc_hd__and2_1 _6958_ (.A(_2926_),
    .B(_2927_),
    .X(_2928_));
 sky130_fd_sc_hd__nor2_1 _6959_ (.A(_2926_),
    .B(_2927_),
    .Y(_2929_));
 sky130_fd_sc_hd__nor2_1 _6960_ (.A(_2928_),
    .B(_2929_),
    .Y(_2930_));
 sky130_fd_sc_hd__xnor2_2 _6961_ (.A(_2887_),
    .B(_2930_),
    .Y(_2931_));
 sky130_fd_sc_hd__a21o_1 _6962_ (.A1(_2819_),
    .A2(_2867_),
    .B1(_2866_),
    .X(_2932_));
 sky130_fd_sc_hd__xor2_2 _6963_ (.A(_2931_),
    .B(_2932_),
    .X(_2933_));
 sky130_fd_sc_hd__xnor2_2 _6964_ (.A(_2817_),
    .B(_2933_),
    .Y(_2934_));
 sky130_fd_sc_hd__or2_1 _6965_ (.A(_2883_),
    .B(_2934_),
    .X(_2935_));
 sky130_fd_sc_hd__and2_1 _6966_ (.A(_2883_),
    .B(_2934_),
    .X(_2936_));
 sky130_fd_sc_hd__xnor2_2 _6967_ (.A(_2883_),
    .B(_2934_),
    .Y(_2937_));
 sky130_fd_sc_hd__a21oi_1 _6968_ (.A1(_2876_),
    .A2(_2878_),
    .B1(_2874_),
    .Y(_2938_));
 sky130_fd_sc_hd__xnor2_2 _6969_ (.A(_2937_),
    .B(_2938_),
    .Y(_2939_));
 sky130_fd_sc_hd__xor2_1 _6970_ (.A(_2882_),
    .B(_2939_),
    .X(\mul_la.reg_p[19] ));
 sky130_fd_sc_hd__a31o_1 _6971_ (.A1(_2061_),
    .A2(_2410_),
    .A3(_2891_),
    .B1(_2894_),
    .X(_2940_));
 sky130_fd_sc_hd__a22o_1 _6972_ (.A1(_2061_),
    .A2(_2487_),
    .B1(_2562_),
    .B2(_2005_),
    .X(_2941_));
 sky130_fd_sc_hd__or4_1 _6973_ (.A(_2006_),
    .B(_2062_),
    .C(_2488_),
    .D(_2563_),
    .X(_2942_));
 sky130_fd_sc_hd__nand2_1 _6974_ (.A(_2941_),
    .B(_2942_),
    .Y(_2943_));
 sky130_fd_sc_hd__nor2_1 _6975_ (.A(net181),
    .B(_2411_),
    .Y(_2944_));
 sky130_fd_sc_hd__or3_1 _6976_ (.A(net181),
    .B(_2411_),
    .C(_2943_),
    .X(_2945_));
 sky130_fd_sc_hd__xnor2_1 _6977_ (.A(_2943_),
    .B(_2944_),
    .Y(_2946_));
 sky130_fd_sc_hd__nand2_1 _6978_ (.A(_2940_),
    .B(_2946_),
    .Y(_2947_));
 sky130_fd_sc_hd__or2_1 _6979_ (.A(_2940_),
    .B(_2946_),
    .X(_2948_));
 sky130_fd_sc_hd__o2bb2a_1 _6980_ (.A1_N(_2947_),
    .A2_N(_2948_),
    .B1(net185),
    .B2(_2644_),
    .X(_2949_));
 sky130_fd_sc_hd__and2b_1 _6981_ (.A_N(_2949_),
    .B(_2899_),
    .X(_2950_));
 sky130_fd_sc_hd__xnor2_1 _6982_ (.A(_2899_),
    .B(_2949_),
    .Y(_2951_));
 sky130_fd_sc_hd__a21o_1 _6983_ (.A1(_2910_),
    .A2(_2919_),
    .B1(_2918_),
    .X(_2952_));
 sky130_fd_sc_hd__a21oi_1 _6984_ (.A1(_2889_),
    .A2(_2897_),
    .B1(_2896_),
    .Y(_2953_));
 sky130_fd_sc_hd__nand2_1 _6985_ (.A(net182),
    .B(_2449_),
    .Y(_2954_));
 sky130_fd_sc_hd__nor2_1 _6986_ (.A(_2142_),
    .B(net178),
    .Y(_2955_));
 sky130_fd_sc_hd__or3_1 _6987_ (.A(net180),
    .B(net178),
    .C(_2954_),
    .X(_2956_));
 sky130_fd_sc_hd__xnor2_1 _6988_ (.A(_2954_),
    .B(_2955_),
    .Y(_2957_));
 sky130_fd_sc_hd__nor2_1 _6989_ (.A(_2025_),
    .B(net225),
    .Y(_2958_));
 sky130_fd_sc_hd__nand2_1 _6990_ (.A(_2957_),
    .B(_2958_),
    .Y(_2959_));
 sky130_fd_sc_hd__xnor2_1 _6991_ (.A(_2957_),
    .B(_2958_),
    .Y(_2960_));
 sky130_fd_sc_hd__o211a_1 _6992_ (.A1(_2260_),
    .A2(_2263_),
    .B1(_1676_),
    .C1(net213),
    .X(_2961_));
 sky130_fd_sc_hd__o211a_1 _6993_ (.A1(_2335_),
    .A2(_2337_),
    .B1(_1680_),
    .C1(net214),
    .X(_2962_));
 sky130_fd_sc_hd__nand2_1 _6994_ (.A(_2961_),
    .B(_2962_),
    .Y(_2963_));
 sky130_fd_sc_hd__xnor2_2 _6995_ (.A(_2961_),
    .B(_2962_),
    .Y(_2964_));
 sky130_fd_sc_hd__nor2_1 _6996_ (.A(_2205_),
    .B(net179),
    .Y(_2965_));
 sky130_fd_sc_hd__xnor2_1 _6997_ (.A(_2964_),
    .B(_2965_),
    .Y(_2966_));
 sky130_fd_sc_hd__o31ai_2 _6998_ (.A1(_2142_),
    .A2(net179),
    .A3(_2914_),
    .B1(_2913_),
    .Y(_2967_));
 sky130_fd_sc_hd__xor2_1 _6999_ (.A(_2966_),
    .B(_2967_),
    .X(_2968_));
 sky130_fd_sc_hd__nand2b_1 _7000_ (.A_N(_2960_),
    .B(_2968_),
    .Y(_2969_));
 sky130_fd_sc_hd__xnor2_1 _7001_ (.A(_2960_),
    .B(_2968_),
    .Y(_2970_));
 sky130_fd_sc_hd__and2b_1 _7002_ (.A_N(_2953_),
    .B(_2970_),
    .X(_2971_));
 sky130_fd_sc_hd__xnor2_1 _7003_ (.A(_2953_),
    .B(_2970_),
    .Y(_2972_));
 sky130_fd_sc_hd__xor2_1 _7004_ (.A(_2952_),
    .B(_2972_),
    .X(_2973_));
 sky130_fd_sc_hd__xnor2_1 _7005_ (.A(_2951_),
    .B(_2973_),
    .Y(_2974_));
 sky130_fd_sc_hd__a21oi_1 _7006_ (.A1(_2901_),
    .A2(_2925_),
    .B1(_2974_),
    .Y(_2975_));
 sky130_fd_sc_hd__and3_1 _7007_ (.A(_2901_),
    .B(_2925_),
    .C(_2974_),
    .X(_2976_));
 sky130_fd_sc_hd__o31a_1 _7008_ (.A1(net168),
    .A2(net225),
    .A3(_2908_),
    .B1(_2907_),
    .X(_2977_));
 sky130_fd_sc_hd__o21bai_1 _7009_ (.A1(_2921_),
    .A2(_2923_),
    .B1_N(_2977_),
    .Y(_2978_));
 sky130_fd_sc_hd__or3b_1 _7010_ (.A(_2921_),
    .B(_2923_),
    .C_N(_2977_),
    .X(_2979_));
 sky130_fd_sc_hd__o2bb2a_1 _7011_ (.A1_N(_2978_),
    .A2_N(_2979_),
    .B1(net168),
    .B2(_2603_),
    .X(_2980_));
 sky130_fd_sc_hd__or3_1 _7012_ (.A(_2975_),
    .B(_2976_),
    .C(_2980_),
    .X(_2981_));
 sky130_fd_sc_hd__o21ai_1 _7013_ (.A1(_2975_),
    .A2(_2976_),
    .B1(_2980_),
    .Y(_2982_));
 sky130_fd_sc_hd__nand2_1 _7014_ (.A(_2981_),
    .B(_2982_),
    .Y(_2983_));
 sky130_fd_sc_hd__o21ba_1 _7015_ (.A1(_2887_),
    .A2(_2929_),
    .B1_N(_2928_),
    .X(_2984_));
 sky130_fd_sc_hd__nor2_1 _7016_ (.A(_2983_),
    .B(_2984_),
    .Y(_2985_));
 sky130_fd_sc_hd__xnor2_1 _7017_ (.A(_2983_),
    .B(_2984_),
    .Y(_2986_));
 sky130_fd_sc_hd__nor2_1 _7018_ (.A(_2885_),
    .B(_2986_),
    .Y(_2987_));
 sky130_fd_sc_hd__and2_1 _7019_ (.A(_2885_),
    .B(_2986_),
    .X(_2988_));
 sky130_fd_sc_hd__nor2_2 _7020_ (.A(_2987_),
    .B(_2988_),
    .Y(_2989_));
 sky130_fd_sc_hd__a32o_2 _7021_ (.A1(_2815_),
    .A2(_2816_),
    .A3(_2933_),
    .B1(_2932_),
    .B2(_2931_),
    .X(_2990_));
 sky130_fd_sc_hd__nand2_1 _7022_ (.A(_2989_),
    .B(_2990_),
    .Y(_2991_));
 sky130_fd_sc_hd__inv_2 _7023_ (.A(_2991_),
    .Y(_2992_));
 sky130_fd_sc_hd__xnor2_2 _7024_ (.A(_2989_),
    .B(_2990_),
    .Y(_2993_));
 sky130_fd_sc_hd__or4_2 _7025_ (.A(_2736_),
    .B(_2811_),
    .C(_2875_),
    .D(_2937_),
    .X(_2994_));
 sky130_fd_sc_hd__a31o_1 _7026_ (.A1(_2737_),
    .A2(_2738_),
    .A3(_2739_),
    .B1(_2994_),
    .X(_2995_));
 sky130_fd_sc_hd__a2111o_1 _7027_ (.A1(_2733_),
    .A2(_2808_),
    .B1(_2809_),
    .C1(_2875_),
    .D1(_2937_),
    .X(_2996_));
 sky130_fd_sc_hd__a21oi_2 _7028_ (.A1(_2874_),
    .A2(_2935_),
    .B1(_2936_),
    .Y(_2997_));
 sky130_fd_sc_hd__and2_1 _7029_ (.A(_2996_),
    .B(_2997_),
    .X(_2998_));
 sky130_fd_sc_hd__a21oi_1 _7030_ (.A1(_2995_),
    .A2(_2998_),
    .B1(_2993_),
    .Y(_2999_));
 sky130_fd_sc_hd__and3_1 _7031_ (.A(_2993_),
    .B(_2995_),
    .C(_2998_),
    .X(_3000_));
 sky130_fd_sc_hd__or2_2 _7032_ (.A(_2999_),
    .B(_3000_),
    .X(_3001_));
 sky130_fd_sc_hd__and4_2 _7033_ (.A(_2742_),
    .B(_2879_),
    .C(_2880_),
    .D(_2939_),
    .X(_3002_));
 sky130_fd_sc_hd__nor2_1 _7034_ (.A(_1809_),
    .B(_3002_),
    .Y(_3003_));
 sky130_fd_sc_hd__xnor2_1 _7035_ (.A(_3001_),
    .B(_3003_),
    .Y(\mul_la.reg_p[20] ));
 sky130_fd_sc_hd__o22a_1 _7036_ (.A1(_2062_),
    .A2(_2563_),
    .B1(_2644_),
    .B2(_2006_),
    .X(_3004_));
 sky130_fd_sc_hd__or3_2 _7037_ (.A(net181),
    .B(_2488_),
    .C(_3004_),
    .X(_3005_));
 sky130_fd_sc_hd__o21ai_1 _7038_ (.A1(net181),
    .A2(_2488_),
    .B1(_3004_),
    .Y(_3006_));
 sky130_fd_sc_hd__and2_1 _7039_ (.A(_3005_),
    .B(_3006_),
    .X(_3007_));
 sky130_fd_sc_hd__nand2_1 _7040_ (.A(_2942_),
    .B(_2945_),
    .Y(_3008_));
 sky130_fd_sc_hd__a21bo_1 _7041_ (.A1(_2942_),
    .A2(_2945_),
    .B1_N(_3007_),
    .X(_3009_));
 sky130_fd_sc_hd__xor2_1 _7042_ (.A(_3007_),
    .B(_3008_),
    .X(_3010_));
 sky130_fd_sc_hd__a21bo_1 _7043_ (.A1(_2966_),
    .A2(_2967_),
    .B1_N(_2969_),
    .X(_3011_));
 sky130_fd_sc_hd__a22o_1 _7044_ (.A1(_2204_),
    .A2(_2376_),
    .B1(_2449_),
    .B2(_2141_),
    .X(_3012_));
 sky130_fd_sc_hd__or4_1 _7045_ (.A(net180),
    .B(_2205_),
    .C(net178),
    .D(_2450_),
    .X(_3013_));
 sky130_fd_sc_hd__nand2_1 _7046_ (.A(_3012_),
    .B(_3013_),
    .Y(_3014_));
 sky130_fd_sc_hd__nand2_1 _7047_ (.A(net182),
    .B(_2523_),
    .Y(_3015_));
 sky130_fd_sc_hd__xor2_1 _7048_ (.A(_3014_),
    .B(_3015_),
    .X(_3016_));
 sky130_fd_sc_hd__o211a_1 _7049_ (.A1(_2335_),
    .A2(_2337_),
    .B1(_1680_),
    .C1(net213),
    .X(_3017_));
 sky130_fd_sc_hd__nand2_1 _7050_ (.A(net214),
    .B(_2410_),
    .Y(_3018_));
 sky130_fd_sc_hd__or3_1 _7051_ (.A(_2235_),
    .B(_2339_),
    .C(_3018_),
    .X(_3019_));
 sky130_fd_sc_hd__xor2_2 _7052_ (.A(_3017_),
    .B(_3018_),
    .X(_3020_));
 sky130_fd_sc_hd__nor2_1 _7053_ (.A(_2265_),
    .B(net179),
    .Y(_3021_));
 sky130_fd_sc_hd__xnor2_1 _7054_ (.A(_3020_),
    .B(_3021_),
    .Y(_3022_));
 sky130_fd_sc_hd__o31ai_2 _7055_ (.A1(_2205_),
    .A2(net179),
    .A3(_2964_),
    .B1(_2963_),
    .Y(_3023_));
 sky130_fd_sc_hd__and2_1 _7056_ (.A(_3022_),
    .B(_3023_),
    .X(_3024_));
 sky130_fd_sc_hd__xor2_1 _7057_ (.A(_3022_),
    .B(_3023_),
    .X(_3025_));
 sky130_fd_sc_hd__xnor2_1 _7058_ (.A(_3016_),
    .B(_3025_),
    .Y(_3026_));
 sky130_fd_sc_hd__nor2_1 _7059_ (.A(_2947_),
    .B(_3026_),
    .Y(_3027_));
 sky130_fd_sc_hd__xnor2_1 _7060_ (.A(_2947_),
    .B(_3026_),
    .Y(_3028_));
 sky130_fd_sc_hd__and2b_1 _7061_ (.A_N(_3028_),
    .B(_3011_),
    .X(_3029_));
 sky130_fd_sc_hd__xnor2_1 _7062_ (.A(_3011_),
    .B(_3028_),
    .Y(_3030_));
 sky130_fd_sc_hd__nand2_1 _7063_ (.A(_3010_),
    .B(_3030_),
    .Y(_3031_));
 sky130_fd_sc_hd__xnor2_1 _7064_ (.A(_3010_),
    .B(_3030_),
    .Y(_3032_));
 sky130_fd_sc_hd__a21oi_1 _7065_ (.A1(_2951_),
    .A2(_2973_),
    .B1(_2950_),
    .Y(_3033_));
 sky130_fd_sc_hd__or2_1 _7066_ (.A(_3032_),
    .B(_3033_),
    .X(_3034_));
 sky130_fd_sc_hd__xnor2_1 _7067_ (.A(_3032_),
    .B(_3033_),
    .Y(_3035_));
 sky130_fd_sc_hd__a21oi_2 _7068_ (.A1(_2952_),
    .A2(_2972_),
    .B1(_2971_),
    .Y(_3036_));
 sky130_fd_sc_hd__a21oi_2 _7069_ (.A1(_2956_),
    .A2(_2959_),
    .B1(_3036_),
    .Y(_3037_));
 sky130_fd_sc_hd__and3_1 _7070_ (.A(_2956_),
    .B(_2959_),
    .C(_3036_),
    .X(_3038_));
 sky130_fd_sc_hd__o22a_1 _7071_ (.A1(_2025_),
    .A2(_2603_),
    .B1(_3037_),
    .B2(_3038_),
    .X(_3039_));
 sky130_fd_sc_hd__xnor2_1 _7072_ (.A(_3035_),
    .B(_3039_),
    .Y(_3040_));
 sky130_fd_sc_hd__o21ba_1 _7073_ (.A1(_2976_),
    .A2(_2980_),
    .B1_N(_2975_),
    .X(_3041_));
 sky130_fd_sc_hd__nor2_1 _7074_ (.A(_3040_),
    .B(_3041_),
    .Y(_3042_));
 sky130_fd_sc_hd__xnor2_1 _7075_ (.A(_3040_),
    .B(_3041_),
    .Y(_3043_));
 sky130_fd_sc_hd__nor2_1 _7076_ (.A(_2978_),
    .B(_3043_),
    .Y(_3044_));
 sky130_fd_sc_hd__and2_1 _7077_ (.A(_2978_),
    .B(_3043_),
    .X(_3045_));
 sky130_fd_sc_hd__nor2_1 _7078_ (.A(_3044_),
    .B(_3045_),
    .Y(_3046_));
 sky130_fd_sc_hd__o21a_1 _7079_ (.A1(_2985_),
    .A2(_2987_),
    .B1(_3046_),
    .X(_3047_));
 sky130_fd_sc_hd__inv_2 _7080_ (.A(_3047_),
    .Y(_3048_));
 sky130_fd_sc_hd__nor3_2 _7081_ (.A(_2985_),
    .B(_2987_),
    .C(_3046_),
    .Y(_3049_));
 sky130_fd_sc_hd__or2_1 _7082_ (.A(_3047_),
    .B(_3049_),
    .X(_3050_));
 sky130_fd_sc_hd__or3_1 _7083_ (.A(_2992_),
    .B(_2999_),
    .C(_3050_),
    .X(_3051_));
 sky130_fd_sc_hd__o21ai_1 _7084_ (.A1(_2992_),
    .A2(_2999_),
    .B1(_3050_),
    .Y(_3052_));
 sky130_fd_sc_hd__and2_1 _7085_ (.A(_3051_),
    .B(_3052_),
    .X(_3053_));
 sky130_fd_sc_hd__a21oi_1 _7086_ (.A1(_3001_),
    .A2(_3002_),
    .B1(_1809_),
    .Y(_3054_));
 sky130_fd_sc_hd__xnor2_1 _7087_ (.A(_3053_),
    .B(_3054_),
    .Y(\mul_la.reg_p[21] ));
 sky130_fd_sc_hd__a22o_1 _7088_ (.A1(_2116_),
    .A2(_2562_),
    .B1(_2643_),
    .B2(_2061_),
    .X(_3055_));
 sky130_fd_sc_hd__and2_1 _7089_ (.A(_3005_),
    .B(_3055_),
    .X(_3056_));
 sky130_fd_sc_hd__a21o_1 _7090_ (.A1(_3016_),
    .A2(_3025_),
    .B1(_3024_),
    .X(_3057_));
 sky130_fd_sc_hd__a22o_1 _7091_ (.A1(_2264_),
    .A2(_2376_),
    .B1(_2449_),
    .B2(_2204_),
    .X(_3058_));
 sky130_fd_sc_hd__or4_1 _7092_ (.A(_2205_),
    .B(_2265_),
    .C(_2377_),
    .D(_2450_),
    .X(_3059_));
 sky130_fd_sc_hd__nand2_1 _7093_ (.A(_3058_),
    .B(_3059_),
    .Y(_3060_));
 sky130_fd_sc_hd__nand2_1 _7094_ (.A(_2141_),
    .B(_2523_),
    .Y(_3061_));
 sky130_fd_sc_hd__xnor2_1 _7095_ (.A(_3060_),
    .B(_3061_),
    .Y(_3062_));
 sky130_fd_sc_hd__a22o_1 _7096_ (.A1(net213),
    .A2(_2410_),
    .B1(_2487_),
    .B2(net214),
    .X(_3063_));
 sky130_fd_sc_hd__nand4_1 _7097_ (.A(net214),
    .B(net213),
    .C(_2410_),
    .D(_2487_),
    .Y(_3064_));
 sky130_fd_sc_hd__nand2_1 _7098_ (.A(_3063_),
    .B(_3064_),
    .Y(_3065_));
 sky130_fd_sc_hd__nand2_1 _7099_ (.A(_2302_),
    .B(_2338_),
    .Y(_3066_));
 sky130_fd_sc_hd__xnor2_1 _7100_ (.A(_3065_),
    .B(_3066_),
    .Y(_3067_));
 sky130_fd_sc_hd__o31ai_2 _7101_ (.A1(_2265_),
    .A2(net179),
    .A3(_3020_),
    .B1(_3019_),
    .Y(_3068_));
 sky130_fd_sc_hd__nand2b_1 _7102_ (.A_N(_3067_),
    .B(_3068_),
    .Y(_3069_));
 sky130_fd_sc_hd__xor2_1 _7103_ (.A(_3067_),
    .B(_3068_),
    .X(_3070_));
 sky130_fd_sc_hd__xnor2_1 _7104_ (.A(_3062_),
    .B(_3070_),
    .Y(_3071_));
 sky130_fd_sc_hd__nor2_1 _7105_ (.A(_3009_),
    .B(_3071_),
    .Y(_3072_));
 sky130_fd_sc_hd__xor2_1 _7106_ (.A(_3009_),
    .B(_3071_),
    .X(_3073_));
 sky130_fd_sc_hd__xor2_1 _7107_ (.A(_3057_),
    .B(_3073_),
    .X(_3074_));
 sky130_fd_sc_hd__nand2_1 _7108_ (.A(_3056_),
    .B(_3074_),
    .Y(_3075_));
 sky130_fd_sc_hd__xnor2_1 _7109_ (.A(_3056_),
    .B(_3074_),
    .Y(_3076_));
 sky130_fd_sc_hd__nor2_1 _7110_ (.A(_3031_),
    .B(_3076_),
    .Y(_3077_));
 sky130_fd_sc_hd__xor2_1 _7111_ (.A(_3031_),
    .B(_3076_),
    .X(_3078_));
 sky130_fd_sc_hd__o21ai_1 _7112_ (.A1(_3014_),
    .A2(_3015_),
    .B1(_3013_),
    .Y(_3079_));
 sky130_fd_sc_hd__o21a_1 _7113_ (.A1(_3027_),
    .A2(_3029_),
    .B1(_3079_),
    .X(_3080_));
 sky130_fd_sc_hd__nor3_1 _7114_ (.A(_3027_),
    .B(_3029_),
    .C(_3079_),
    .Y(_3081_));
 sky130_fd_sc_hd__a2bb2o_1 _7115_ (.A1_N(_3080_),
    .A2_N(_3081_),
    .B1(net182),
    .B2(_2602_),
    .X(_3082_));
 sky130_fd_sc_hd__and2_1 _7116_ (.A(_3078_),
    .B(_3082_),
    .X(_3083_));
 sky130_fd_sc_hd__nor2_1 _7117_ (.A(_3078_),
    .B(_3082_),
    .Y(_3084_));
 sky130_fd_sc_hd__nor2_1 _7118_ (.A(_3083_),
    .B(_3084_),
    .Y(_3085_));
 sky130_fd_sc_hd__o21a_1 _7119_ (.A1(_3035_),
    .A2(_3039_),
    .B1(_3034_),
    .X(_3086_));
 sky130_fd_sc_hd__or3_1 _7120_ (.A(_3083_),
    .B(_3084_),
    .C(_3086_),
    .X(_3087_));
 sky130_fd_sc_hd__xnor2_1 _7121_ (.A(_3085_),
    .B(_3086_),
    .Y(_3088_));
 sky130_fd_sc_hd__nand2_1 _7122_ (.A(_3037_),
    .B(_3088_),
    .Y(_3089_));
 sky130_fd_sc_hd__xor2_1 _7123_ (.A(_3037_),
    .B(_3088_),
    .X(_3090_));
 sky130_fd_sc_hd__o21ai_2 _7124_ (.A1(_3042_),
    .A2(_3044_),
    .B1(_3090_),
    .Y(_3091_));
 sky130_fd_sc_hd__or3_1 _7125_ (.A(_3042_),
    .B(_3044_),
    .C(_3090_),
    .X(_3092_));
 sky130_fd_sc_hd__nand2_2 _7126_ (.A(_3091_),
    .B(_3092_),
    .Y(_3093_));
 sky130_fd_sc_hd__a21o_1 _7127_ (.A1(_2991_),
    .A2(_3048_),
    .B1(_3049_),
    .X(_3094_));
 sky130_fd_sc_hd__a21o_1 _7128_ (.A1(_2995_),
    .A2(_2998_),
    .B1(_3050_),
    .X(_3095_));
 sky130_fd_sc_hd__o21a_1 _7129_ (.A1(_2993_),
    .A2(_3095_),
    .B1(_3094_),
    .X(_3096_));
 sky130_fd_sc_hd__xor2_2 _7130_ (.A(_3093_),
    .B(_3096_),
    .X(_3097_));
 sky130_fd_sc_hd__nand3_1 _7131_ (.A(_3001_),
    .B(_3051_),
    .C(_3052_),
    .Y(_3098_));
 sky130_fd_sc_hd__a31o_1 _7132_ (.A1(_3001_),
    .A2(_3002_),
    .A3(_3053_),
    .B1(_1809_),
    .X(_3099_));
 sky130_fd_sc_hd__xnor2_1 _7133_ (.A(_3097_),
    .B(_3099_),
    .Y(\mul_la.reg_p[22] ));
 sky130_fd_sc_hd__nor2_1 _7134_ (.A(_3097_),
    .B(_3098_),
    .Y(_3100_));
 sky130_fd_sc_hd__a21oi_1 _7135_ (.A1(_3002_),
    .A2(_3100_),
    .B1(_1809_),
    .Y(_3101_));
 sky130_fd_sc_hd__o21ai_1 _7136_ (.A1(_3062_),
    .A2(_3070_),
    .B1(_3069_),
    .Y(_3102_));
 sky130_fd_sc_hd__a22o_1 _7137_ (.A1(_2338_),
    .A2(_2376_),
    .B1(_2449_),
    .B2(_2264_),
    .X(_3103_));
 sky130_fd_sc_hd__or4_1 _7138_ (.A(_2265_),
    .B(_2339_),
    .C(_2377_),
    .D(_2450_),
    .X(_3104_));
 sky130_fd_sc_hd__nand2_1 _7139_ (.A(_3103_),
    .B(_3104_),
    .Y(_3105_));
 sky130_fd_sc_hd__nor2_1 _7140_ (.A(_2205_),
    .B(net225),
    .Y(_3106_));
 sky130_fd_sc_hd__xnor2_2 _7141_ (.A(_3105_),
    .B(_3106_),
    .Y(_3107_));
 sky130_fd_sc_hd__a22oi_2 _7142_ (.A1(net213),
    .A2(_2487_),
    .B1(_2562_),
    .B2(net214),
    .Y(_3108_));
 sky130_fd_sc_hd__and4_1 _7143_ (.A(net214),
    .B(net213),
    .C(_2487_),
    .D(_2562_),
    .X(_3109_));
 sky130_fd_sc_hd__nor2_1 _7144_ (.A(_3108_),
    .B(_3109_),
    .Y(_3110_));
 sky130_fd_sc_hd__nand2_1 _7145_ (.A(_2302_),
    .B(_2410_),
    .Y(_3111_));
 sky130_fd_sc_hd__xor2_1 _7146_ (.A(_3110_),
    .B(_3111_),
    .X(_3112_));
 sky130_fd_sc_hd__o21ai_1 _7147_ (.A1(_3065_),
    .A2(_3066_),
    .B1(_3064_),
    .Y(_3113_));
 sky130_fd_sc_hd__and2b_1 _7148_ (.A_N(_3112_),
    .B(_3113_),
    .X(_3114_));
 sky130_fd_sc_hd__xnor2_1 _7149_ (.A(_3112_),
    .B(_3113_),
    .Y(_3115_));
 sky130_fd_sc_hd__and2_1 _7150_ (.A(_3107_),
    .B(_3115_),
    .X(_3116_));
 sky130_fd_sc_hd__nor2_1 _7151_ (.A(_3107_),
    .B(_3115_),
    .Y(_3117_));
 sky130_fd_sc_hd__xor2_1 _7152_ (.A(_3107_),
    .B(_3115_),
    .X(_3118_));
 sky130_fd_sc_hd__xnor2_1 _7153_ (.A(_3005_),
    .B(_3118_),
    .Y(_3119_));
 sky130_fd_sc_hd__nand2_1 _7154_ (.A(_3102_),
    .B(_3119_),
    .Y(_3120_));
 sky130_fd_sc_hd__or2_1 _7155_ (.A(_3102_),
    .B(_3119_),
    .X(_3121_));
 sky130_fd_sc_hd__o2bb2a_1 _7156_ (.A1_N(_3120_),
    .A2_N(_3121_),
    .B1(net181),
    .B2(_2644_),
    .X(_3122_));
 sky130_fd_sc_hd__or2_1 _7157_ (.A(_3075_),
    .B(_3122_),
    .X(_3123_));
 sky130_fd_sc_hd__xnor2_1 _7158_ (.A(_3075_),
    .B(_3122_),
    .Y(_3124_));
 sky130_fd_sc_hd__a21oi_1 _7159_ (.A1(_3057_),
    .A2(_3073_),
    .B1(_3072_),
    .Y(_3125_));
 sky130_fd_sc_hd__o31a_1 _7160_ (.A1(net180),
    .A2(net225),
    .A3(_3060_),
    .B1(_3059_),
    .X(_3126_));
 sky130_fd_sc_hd__nor2_1 _7161_ (.A(_3125_),
    .B(_3126_),
    .Y(_3127_));
 sky130_fd_sc_hd__xnor2_1 _7162_ (.A(_3125_),
    .B(_3126_),
    .Y(_3128_));
 sky130_fd_sc_hd__o21a_1 _7163_ (.A1(net180),
    .A2(_2603_),
    .B1(_3128_),
    .X(_3129_));
 sky130_fd_sc_hd__xor2_1 _7164_ (.A(_3124_),
    .B(_3129_),
    .X(_3130_));
 sky130_fd_sc_hd__o21a_1 _7165_ (.A1(_3077_),
    .A2(_3083_),
    .B1(_3130_),
    .X(_3131_));
 sky130_fd_sc_hd__nor3_1 _7166_ (.A(_3077_),
    .B(_3083_),
    .C(_3130_),
    .Y(_3132_));
 sky130_fd_sc_hd__nor2_1 _7167_ (.A(_3131_),
    .B(_3132_),
    .Y(_3133_));
 sky130_fd_sc_hd__xnor2_1 _7168_ (.A(_3080_),
    .B(_3133_),
    .Y(_3134_));
 sky130_fd_sc_hd__nand3_2 _7169_ (.A(_3087_),
    .B(_3089_),
    .C(_3134_),
    .Y(_3135_));
 sky130_fd_sc_hd__a21o_1 _7170_ (.A1(_3087_),
    .A2(_3089_),
    .B1(_3134_),
    .X(_3136_));
 sky130_fd_sc_hd__nand2_2 _7171_ (.A(_3135_),
    .B(_3136_),
    .Y(_3137_));
 sky130_fd_sc_hd__o21ai_2 _7172_ (.A1(_3093_),
    .A2(_3096_),
    .B1(_3091_),
    .Y(_3138_));
 sky130_fd_sc_hd__xor2_4 _7173_ (.A(_3137_),
    .B(_3138_),
    .X(_3139_));
 sky130_fd_sc_hd__xnor2_1 _7174_ (.A(_3101_),
    .B(_3139_),
    .Y(\mul_la.reg_p[23] ));
 sky130_fd_sc_hd__a22o_1 _7175_ (.A1(_2376_),
    .A2(_2410_),
    .B1(_2449_),
    .B2(_2338_),
    .X(_3140_));
 sky130_fd_sc_hd__or4_1 _7176_ (.A(_2339_),
    .B(net178),
    .C(_2411_),
    .D(_2450_),
    .X(_3141_));
 sky130_fd_sc_hd__nand2_1 _7177_ (.A(_3140_),
    .B(_3141_),
    .Y(_3142_));
 sky130_fd_sc_hd__nor2_1 _7178_ (.A(_2265_),
    .B(net225),
    .Y(_3143_));
 sky130_fd_sc_hd__xnor2_1 _7179_ (.A(_3142_),
    .B(_3143_),
    .Y(_3144_));
 sky130_fd_sc_hd__o22a_1 _7180_ (.A1(_2235_),
    .A2(_2563_),
    .B1(_2644_),
    .B2(_2176_),
    .X(_3145_));
 sky130_fd_sc_hd__or3_1 _7181_ (.A(net179),
    .B(_2488_),
    .C(_3145_),
    .X(_3146_));
 sky130_fd_sc_hd__o21ai_1 _7182_ (.A1(net179),
    .A2(_2488_),
    .B1(_3145_),
    .Y(_3147_));
 sky130_fd_sc_hd__and2_1 _7183_ (.A(_3146_),
    .B(_3147_),
    .X(_3148_));
 sky130_fd_sc_hd__o21ba_1 _7184_ (.A1(_3108_),
    .A2(_3111_),
    .B1_N(_3109_),
    .X(_3149_));
 sky130_fd_sc_hd__nand2b_1 _7185_ (.A_N(_3149_),
    .B(_3148_),
    .Y(_3150_));
 sky130_fd_sc_hd__xnor2_1 _7186_ (.A(_3148_),
    .B(_3149_),
    .Y(_3151_));
 sky130_fd_sc_hd__nand2_1 _7187_ (.A(_3144_),
    .B(_3151_),
    .Y(_3152_));
 sky130_fd_sc_hd__or2_1 _7188_ (.A(_3144_),
    .B(_3151_),
    .X(_3153_));
 sky130_fd_sc_hd__nand2_1 _7189_ (.A(_3152_),
    .B(_3153_),
    .Y(_3154_));
 sky130_fd_sc_hd__o211a_1 _7190_ (.A1(_3114_),
    .A2(_3116_),
    .B1(_3152_),
    .C1(_3153_),
    .X(_3155_));
 sky130_fd_sc_hd__or3b_1 _7191_ (.A(_3114_),
    .B(_3116_),
    .C_N(_3154_),
    .X(_3156_));
 sky130_fd_sc_hd__nand2b_1 _7192_ (.A_N(_3155_),
    .B(_3156_),
    .Y(_3157_));
 sky130_fd_sc_hd__o31a_1 _7193_ (.A1(_3005_),
    .A2(_3116_),
    .A3(_3117_),
    .B1(_3120_),
    .X(_3158_));
 sky130_fd_sc_hd__o31a_1 _7194_ (.A1(_2205_),
    .A2(net225),
    .A3(_3105_),
    .B1(_3104_),
    .X(_3159_));
 sky130_fd_sc_hd__or2_1 _7195_ (.A(_3158_),
    .B(_3159_),
    .X(_3160_));
 sky130_fd_sc_hd__xnor2_1 _7196_ (.A(_3158_),
    .B(_3159_),
    .Y(_3161_));
 sky130_fd_sc_hd__nand2_1 _7197_ (.A(_2204_),
    .B(_2602_),
    .Y(_3162_));
 sky130_fd_sc_hd__a21o_1 _7198_ (.A1(_3161_),
    .A2(_3162_),
    .B1(_3157_),
    .X(_3163_));
 sky130_fd_sc_hd__nand3_1 _7199_ (.A(_3157_),
    .B(_3161_),
    .C(_3162_),
    .Y(_3164_));
 sky130_fd_sc_hd__nand2_1 _7200_ (.A(_3163_),
    .B(_3164_),
    .Y(_3165_));
 sky130_fd_sc_hd__o21a_1 _7201_ (.A1(_3124_),
    .A2(_3129_),
    .B1(_3123_),
    .X(_3166_));
 sky130_fd_sc_hd__nor2_1 _7202_ (.A(_3165_),
    .B(_3166_),
    .Y(_3167_));
 sky130_fd_sc_hd__xor2_1 _7203_ (.A(_3165_),
    .B(_3166_),
    .X(_3168_));
 sky130_fd_sc_hd__and2_1 _7204_ (.A(_3127_),
    .B(_3168_),
    .X(_3169_));
 sky130_fd_sc_hd__nor2_1 _7205_ (.A(_3127_),
    .B(_3168_),
    .Y(_3170_));
 sky130_fd_sc_hd__nor2_1 _7206_ (.A(_3169_),
    .B(_3170_),
    .Y(_3171_));
 sky130_fd_sc_hd__a21o_1 _7207_ (.A1(_3080_),
    .A2(_3133_),
    .B1(_3131_),
    .X(_3172_));
 sky130_fd_sc_hd__nand2_1 _7208_ (.A(_3171_),
    .B(_3172_),
    .Y(_3173_));
 sky130_fd_sc_hd__or2_1 _7209_ (.A(_3171_),
    .B(_3172_),
    .X(_3174_));
 sky130_fd_sc_hd__and2_1 _7210_ (.A(_3173_),
    .B(_3174_),
    .X(_3175_));
 sky130_fd_sc_hd__or4_1 _7211_ (.A(_2993_),
    .B(_3050_),
    .C(_3093_),
    .D(_3137_),
    .X(_3176_));
 sky130_fd_sc_hd__a21o_1 _7212_ (.A1(_2996_),
    .A2(_2997_),
    .B1(_3176_),
    .X(_3177_));
 sky130_fd_sc_hd__a311o_1 _7213_ (.A1(_2737_),
    .A2(_2738_),
    .A3(_2739_),
    .B1(_2994_),
    .C1(_3176_),
    .X(_3178_));
 sky130_fd_sc_hd__nand2b_1 _7214_ (.A_N(_3091_),
    .B(_3135_),
    .Y(_3179_));
 sky130_fd_sc_hd__o311a_1 _7215_ (.A1(_3093_),
    .A2(_3094_),
    .A3(_3137_),
    .B1(_3179_),
    .C1(_3136_),
    .X(_3180_));
 sky130_fd_sc_hd__nand3_2 _7216_ (.A(_3177_),
    .B(_3178_),
    .C(_3180_),
    .Y(_3181_));
 sky130_fd_sc_hd__xor2_2 _7217_ (.A(_3175_),
    .B(_3181_),
    .X(_3182_));
 sky130_fd_sc_hd__nand3_2 _7218_ (.A(_3002_),
    .B(_3100_),
    .C(_3139_),
    .Y(_3183_));
 sky130_fd_sc_hd__nand2_1 _7219_ (.A(net251),
    .B(_3183_),
    .Y(_3184_));
 sky130_fd_sc_hd__xnor2_1 _7220_ (.A(_3182_),
    .B(_3184_),
    .Y(\mul_la.reg_p[24] ));
 sky130_fd_sc_hd__o22a_1 _7221_ (.A1(_2411_),
    .A2(_2450_),
    .B1(_2488_),
    .B2(net178),
    .X(_3185_));
 sky130_fd_sc_hd__and4_1 _7222_ (.A(_2376_),
    .B(_2410_),
    .C(_2449_),
    .D(_2487_),
    .X(_3186_));
 sky130_fd_sc_hd__nor2_1 _7223_ (.A(_3185_),
    .B(_3186_),
    .Y(_3187_));
 sky130_fd_sc_hd__nor2_1 _7224_ (.A(_2339_),
    .B(net225),
    .Y(_3188_));
 sky130_fd_sc_hd__xnor2_1 _7225_ (.A(_3187_),
    .B(_3188_),
    .Y(_3189_));
 sky130_fd_sc_hd__a22o_1 _7226_ (.A1(_2302_),
    .A2(_2562_),
    .B1(_2643_),
    .B2(net213),
    .X(_3190_));
 sky130_fd_sc_hd__nand2_1 _7227_ (.A(_3146_),
    .B(_3190_),
    .Y(_3191_));
 sky130_fd_sc_hd__or2_1 _7228_ (.A(_3189_),
    .B(_3191_),
    .X(_3192_));
 sky130_fd_sc_hd__nand2_1 _7229_ (.A(_3189_),
    .B(_3191_),
    .Y(_3193_));
 sky130_fd_sc_hd__nand2_1 _7230_ (.A(_3192_),
    .B(_3193_),
    .Y(_3194_));
 sky130_fd_sc_hd__a21o_1 _7231_ (.A1(_3150_),
    .A2(_3152_),
    .B1(_3194_),
    .X(_3195_));
 sky130_fd_sc_hd__nand3_1 _7232_ (.A(_3150_),
    .B(_3152_),
    .C(_3194_),
    .Y(_3196_));
 sky130_fd_sc_hd__and2_1 _7233_ (.A(_3195_),
    .B(_3196_),
    .X(_3197_));
 sky130_fd_sc_hd__a21bo_1 _7234_ (.A1(_3140_),
    .A2(_3143_),
    .B1_N(_3141_),
    .X(_3198_));
 sky130_fd_sc_hd__nand2_1 _7235_ (.A(_3155_),
    .B(_3198_),
    .Y(_3199_));
 sky130_fd_sc_hd__xor2_1 _7236_ (.A(_3155_),
    .B(_3198_),
    .X(_3200_));
 sky130_fd_sc_hd__nor2_1 _7237_ (.A(_2265_),
    .B(_2603_),
    .Y(_3201_));
 sky130_fd_sc_hd__o21ai_1 _7238_ (.A1(_3200_),
    .A2(_3201_),
    .B1(_3197_),
    .Y(_3202_));
 sky130_fd_sc_hd__or3_1 _7239_ (.A(_3197_),
    .B(_3200_),
    .C(_3201_),
    .X(_3203_));
 sky130_fd_sc_hd__and2_1 _7240_ (.A(_3202_),
    .B(_3203_),
    .X(_3204_));
 sky130_fd_sc_hd__and2b_1 _7241_ (.A_N(_3163_),
    .B(_3204_),
    .X(_3205_));
 sky130_fd_sc_hd__xnor2_1 _7242_ (.A(_3163_),
    .B(_3204_),
    .Y(_3206_));
 sky130_fd_sc_hd__and2b_1 _7243_ (.A_N(_3160_),
    .B(_3206_),
    .X(_3207_));
 sky130_fd_sc_hd__xnor2_1 _7244_ (.A(_3160_),
    .B(_3206_),
    .Y(_3208_));
 sky130_fd_sc_hd__o21ai_2 _7245_ (.A1(_3167_),
    .A2(_3169_),
    .B1(_3208_),
    .Y(_3209_));
 sky130_fd_sc_hd__or3_1 _7246_ (.A(_3167_),
    .B(_3169_),
    .C(_3208_),
    .X(_3210_));
 sky130_fd_sc_hd__and2_1 _7247_ (.A(_3209_),
    .B(_3210_),
    .X(_3211_));
 sky130_fd_sc_hd__a21bo_1 _7248_ (.A1(_3175_),
    .A2(_3181_),
    .B1_N(_3173_),
    .X(_3212_));
 sky130_fd_sc_hd__xor2_2 _7249_ (.A(_3211_),
    .B(_3212_),
    .X(_3213_));
 sky130_fd_sc_hd__o21ai_1 _7250_ (.A1(_3182_),
    .A2(_3183_),
    .B1(net251),
    .Y(_3214_));
 sky130_fd_sc_hd__xnor2_1 _7251_ (.A(_3213_),
    .B(_3214_),
    .Y(\mul_la.reg_p[25] ));
 sky130_fd_sc_hd__o22a_1 _7252_ (.A1(_2450_),
    .A2(_2488_),
    .B1(_2563_),
    .B2(net178),
    .X(_3215_));
 sky130_fd_sc_hd__or4_1 _7253_ (.A(net178),
    .B(_2450_),
    .C(_2488_),
    .D(_2563_),
    .X(_3216_));
 sky130_fd_sc_hd__and2b_1 _7254_ (.A_N(_3215_),
    .B(_3216_),
    .X(_3217_));
 sky130_fd_sc_hd__nor2_1 _7255_ (.A(_2411_),
    .B(net225),
    .Y(_3218_));
 sky130_fd_sc_hd__xnor2_1 _7256_ (.A(_3217_),
    .B(_3218_),
    .Y(_3219_));
 sky130_fd_sc_hd__o21a_1 _7257_ (.A1(net179),
    .A2(_2644_),
    .B1(_3219_),
    .X(_3220_));
 sky130_fd_sc_hd__a21oi_1 _7258_ (.A1(_3146_),
    .A2(_3192_),
    .B1(_3220_),
    .Y(_3221_));
 sky130_fd_sc_hd__and3_1 _7259_ (.A(_3146_),
    .B(_3192_),
    .C(_3220_),
    .X(_3222_));
 sky130_fd_sc_hd__or2_1 _7260_ (.A(_3221_),
    .B(_3222_),
    .X(_3223_));
 sky130_fd_sc_hd__a21oi_1 _7261_ (.A1(_3187_),
    .A2(_3188_),
    .B1(_3186_),
    .Y(_3224_));
 sky130_fd_sc_hd__nor2_1 _7262_ (.A(_3195_),
    .B(_3224_),
    .Y(_3225_));
 sky130_fd_sc_hd__inv_2 _7263_ (.A(_3225_),
    .Y(_3226_));
 sky130_fd_sc_hd__nand2_1 _7264_ (.A(_3195_),
    .B(_3224_),
    .Y(_3227_));
 sky130_fd_sc_hd__o2bb2a_1 _7265_ (.A1_N(_3226_),
    .A2_N(_3227_),
    .B1(_2339_),
    .B2(_2603_),
    .X(_3228_));
 sky130_fd_sc_hd__nor2_1 _7266_ (.A(_3223_),
    .B(_3228_),
    .Y(_3229_));
 sky130_fd_sc_hd__and2_1 _7267_ (.A(_3223_),
    .B(_3228_),
    .X(_3230_));
 sky130_fd_sc_hd__or2_1 _7268_ (.A(_3229_),
    .B(_3230_),
    .X(_3231_));
 sky130_fd_sc_hd__nor2_1 _7269_ (.A(_3202_),
    .B(_3231_),
    .Y(_3232_));
 sky130_fd_sc_hd__and2_1 _7270_ (.A(_3202_),
    .B(_3231_),
    .X(_3233_));
 sky130_fd_sc_hd__or2_1 _7271_ (.A(_3232_),
    .B(_3233_),
    .X(_3234_));
 sky130_fd_sc_hd__nor2_1 _7272_ (.A(_3199_),
    .B(_3234_),
    .Y(_3235_));
 sky130_fd_sc_hd__and2_1 _7273_ (.A(_3199_),
    .B(_3234_),
    .X(_3236_));
 sky130_fd_sc_hd__nor2_1 _7274_ (.A(_3235_),
    .B(_3236_),
    .Y(_3237_));
 sky130_fd_sc_hd__or2_1 _7275_ (.A(_3205_),
    .B(_3207_),
    .X(_3238_));
 sky130_fd_sc_hd__nand2_1 _7276_ (.A(_3237_),
    .B(_3238_),
    .Y(_3239_));
 sky130_fd_sc_hd__or2_1 _7277_ (.A(_3237_),
    .B(_3238_),
    .X(_3240_));
 sky130_fd_sc_hd__nand2_1 _7278_ (.A(_3239_),
    .B(_3240_),
    .Y(_3241_));
 sky130_fd_sc_hd__nand2_1 _7279_ (.A(_3175_),
    .B(_3211_),
    .Y(_3242_));
 sky130_fd_sc_hd__a31o_1 _7280_ (.A1(_3177_),
    .A2(_3178_),
    .A3(_3180_),
    .B1(_3242_),
    .X(_3243_));
 sky130_fd_sc_hd__a21bo_1 _7281_ (.A1(_3173_),
    .A2(_3209_),
    .B1_N(_3210_),
    .X(_3244_));
 sky130_fd_sc_hd__a21o_2 _7282_ (.A1(_3243_),
    .A2(_3244_),
    .B1(_3241_),
    .X(_3245_));
 sky130_fd_sc_hd__nand3_1 _7283_ (.A(_3241_),
    .B(_3243_),
    .C(_3244_),
    .Y(_3246_));
 sky130_fd_sc_hd__and2_1 _7284_ (.A(_3245_),
    .B(_3246_),
    .X(_3247_));
 sky130_fd_sc_hd__o31ai_1 _7285_ (.A1(_3182_),
    .A2(_3183_),
    .A3(_3213_),
    .B1(net251),
    .Y(_3248_));
 sky130_fd_sc_hd__xnor2_1 _7286_ (.A(_3247_),
    .B(_3248_),
    .Y(\mul_la.reg_p[26] ));
 sky130_fd_sc_hd__a21bo_1 _7287_ (.A1(_3217_),
    .A2(_3218_),
    .B1_N(_3216_),
    .X(_3249_));
 sky130_fd_sc_hd__nand2_1 _7288_ (.A(_3221_),
    .B(_3249_),
    .Y(_3250_));
 sky130_fd_sc_hd__or2_1 _7289_ (.A(_3221_),
    .B(_3249_),
    .X(_3251_));
 sky130_fd_sc_hd__and2_1 _7290_ (.A(_3250_),
    .B(_3251_),
    .X(_3252_));
 sky130_fd_sc_hd__nor2_1 _7291_ (.A(_2411_),
    .B(_2603_),
    .Y(_3253_));
 sky130_fd_sc_hd__o22a_1 _7292_ (.A1(_2450_),
    .A2(_2563_),
    .B1(_2644_),
    .B2(net178),
    .X(_3254_));
 sky130_fd_sc_hd__o21a_1 _7293_ (.A1(_2488_),
    .A2(net225),
    .B1(_3254_),
    .X(_3255_));
 sky130_fd_sc_hd__and3b_1 _7294_ (.A_N(_3254_),
    .B(_2523_),
    .C(_2487_),
    .X(_3256_));
 sky130_fd_sc_hd__nor2_1 _7295_ (.A(_3255_),
    .B(_3256_),
    .Y(_3257_));
 sky130_fd_sc_hd__o21a_1 _7296_ (.A1(_3252_),
    .A2(_3253_),
    .B1(_3257_),
    .X(_3258_));
 sky130_fd_sc_hd__or3_1 _7297_ (.A(_3252_),
    .B(_3253_),
    .C(_3257_),
    .X(_3259_));
 sky130_fd_sc_hd__and2b_1 _7298_ (.A_N(_3258_),
    .B(_3259_),
    .X(_3260_));
 sky130_fd_sc_hd__nand2_1 _7299_ (.A(_3229_),
    .B(_3260_),
    .Y(_3261_));
 sky130_fd_sc_hd__or2_1 _7300_ (.A(_3229_),
    .B(_3260_),
    .X(_3262_));
 sky130_fd_sc_hd__nand2_1 _7301_ (.A(_3261_),
    .B(_3262_),
    .Y(_3263_));
 sky130_fd_sc_hd__xnor2_1 _7302_ (.A(_3225_),
    .B(_3263_),
    .Y(_3264_));
 sky130_fd_sc_hd__or3_1 _7303_ (.A(_3232_),
    .B(_3235_),
    .C(_3264_),
    .X(_3265_));
 sky130_fd_sc_hd__inv_2 _7304_ (.A(_3265_),
    .Y(_3266_));
 sky130_fd_sc_hd__o21a_1 _7305_ (.A1(_3232_),
    .A2(_3235_),
    .B1(_3264_),
    .X(_3267_));
 sky130_fd_sc_hd__nor2_1 _7306_ (.A(_3266_),
    .B(_3267_),
    .Y(_3268_));
 sky130_fd_sc_hd__inv_2 _7307_ (.A(_3268_),
    .Y(_3269_));
 sky130_fd_sc_hd__nand2_1 _7308_ (.A(_3239_),
    .B(_3245_),
    .Y(_3270_));
 sky130_fd_sc_hd__xnor2_2 _7309_ (.A(_3268_),
    .B(_3270_),
    .Y(_3271_));
 sky130_fd_sc_hd__or3_2 _7310_ (.A(_3182_),
    .B(_3213_),
    .C(_3247_),
    .X(_3272_));
 sky130_fd_sc_hd__o21a_1 _7311_ (.A1(_3183_),
    .A2(_3272_),
    .B1(net700),
    .X(_3273_));
 sky130_fd_sc_hd__xnor2_1 _7312_ (.A(_3271_),
    .B(_3273_),
    .Y(\mul_la.reg_p[27] ));
 sky130_fd_sc_hd__nand2_1 _7313_ (.A(net236),
    .B(_2562_),
    .Y(_3274_));
 sky130_fd_sc_hd__o221a_1 _7314_ (.A1(_2488_),
    .A2(_2603_),
    .B1(_2644_),
    .B2(_2450_),
    .C1(_3274_),
    .X(_3275_));
 sky130_fd_sc_hd__nor2_1 _7315_ (.A(_3256_),
    .B(_3275_),
    .Y(_3276_));
 sky130_fd_sc_hd__xnor2_1 _7316_ (.A(_3258_),
    .B(_3276_),
    .Y(_3277_));
 sky130_fd_sc_hd__o21a_1 _7317_ (.A1(_3226_),
    .A2(_3263_),
    .B1(_3261_),
    .X(_3278_));
 sky130_fd_sc_hd__a21o_1 _7318_ (.A1(_3250_),
    .A2(_3277_),
    .B1(_3278_),
    .X(_3279_));
 sky130_fd_sc_hd__nand3_1 _7319_ (.A(_3250_),
    .B(_3277_),
    .C(_3278_),
    .Y(_3280_));
 sky130_fd_sc_hd__nand2_2 _7320_ (.A(_3279_),
    .B(_3280_),
    .Y(_3281_));
 sky130_fd_sc_hd__o21ba_1 _7321_ (.A1(_3239_),
    .A2(_3266_),
    .B1_N(_3267_),
    .X(_3282_));
 sky130_fd_sc_hd__o21ai_4 _7322_ (.A1(_3245_),
    .A2(_3269_),
    .B1(_3282_),
    .Y(_3283_));
 sky130_fd_sc_hd__nand2b_1 _7323_ (.A_N(_3281_),
    .B(_3283_),
    .Y(_3284_));
 sky130_fd_sc_hd__xor2_4 _7324_ (.A(_3281_),
    .B(_3283_),
    .X(_3285_));
 sky130_fd_sc_hd__inv_2 _7325_ (.A(_3285_),
    .Y(_3286_));
 sky130_fd_sc_hd__nand4_2 _7326_ (.A(_3002_),
    .B(_3100_),
    .C(_3139_),
    .D(_3271_),
    .Y(_3287_));
 sky130_fd_sc_hd__o21a_1 _7327_ (.A1(_3272_),
    .A2(_3287_),
    .B1(net700),
    .X(_3288_));
 sky130_fd_sc_hd__xnor2_1 _7328_ (.A(_3285_),
    .B(_3288_),
    .Y(\mul_la.reg_p[28] ));
 sky130_fd_sc_hd__a221o_1 _7329_ (.A1(_1693_),
    .A2(_2602_),
    .B1(_2643_),
    .B2(net236),
    .C1(_3256_),
    .X(_3289_));
 sky130_fd_sc_hd__a21oi_1 _7330_ (.A1(_3258_),
    .A2(_3276_),
    .B1(_3289_),
    .Y(_3290_));
 sky130_fd_sc_hd__and3_1 _7331_ (.A(_3279_),
    .B(_3284_),
    .C(_3290_),
    .X(_3291_));
 sky130_fd_sc_hd__o31a_1 _7332_ (.A1(_3272_),
    .A2(_3286_),
    .A3(_3287_),
    .B1(net251),
    .X(_3292_));
 sky130_fd_sc_hd__xnor2_1 _7333_ (.A(_3291_),
    .B(_3292_),
    .Y(\mul_la.reg_p[29] ));
 sky130_fd_sc_hd__and4_1 _7334_ (.A(_3279_),
    .B(_3284_),
    .C(_3285_),
    .D(_3290_),
    .X(_3293_));
 sky130_fd_sc_hd__or3b_4 _7335_ (.A(_3272_),
    .B(_3287_),
    .C_N(_3293_),
    .X(_3294_));
 sky130_fd_sc_hd__and2_1 _7336_ (.A(net251),
    .B(_3294_),
    .X(\mul_la.reg_p[31] ));
 sky130_fd_sc_hd__a32o_1 _7337_ (.A1(_1572_),
    .A2(_1574_),
    .A3(_2643_),
    .B1(_3294_),
    .B2(net251),
    .X(\mul_la.reg_p[30] ));
 sky130_fd_sc_hd__or4bb_1 _7338_ (.A(net74),
    .B(net73),
    .C_N(net70),
    .D_N(net71),
    .X(_3295_));
 sky130_fd_sc_hd__or4_1 _7339_ (.A(net67),
    .B(net66),
    .C(net69),
    .D(net427),
    .X(_3296_));
 sky130_fd_sc_hd__or4_1 _7340_ (.A(net63),
    .B(net62),
    .C(net65),
    .D(net64),
    .X(_3297_));
 sky130_fd_sc_hd__or4_1 _7341_ (.A(net81),
    .B(net80),
    .C(net52),
    .D(net51),
    .X(_3298_));
 sky130_fd_sc_hd__or4_1 _7342_ (.A(net77),
    .B(net76),
    .C(net79),
    .D(net78),
    .X(_3299_));
 sky130_fd_sc_hd__or4_1 _7343_ (.A(net54),
    .B(net53),
    .C(net56),
    .D(net55),
    .X(_3300_));
 sky130_fd_sc_hd__or4_1 _7344_ (.A(net58),
    .B(net57),
    .C(net60),
    .D(net59),
    .X(_3301_));
 sky130_fd_sc_hd__or4_1 _7345_ (.A(_3298_),
    .B(_3299_),
    .C(_3300_),
    .D(_3301_),
    .X(_3302_));
 sky130_fd_sc_hd__nor4_1 _7346_ (.A(_3295_),
    .B(net428),
    .C(net967),
    .D(_3302_),
    .Y(_3303_));
 sky130_fd_sc_hd__nor2_1 _7347_ (.A(net392),
    .B(net50),
    .Y(_3304_));
 sky130_fd_sc_hd__and4_1 _7348_ (.A(net99),
    .B(net278),
    .C(net429),
    .D(net393),
    .X(_0160_));
 sky130_fd_sc_hd__nand2_1 _7349_ (.A(net396),
    .B(net429),
    .Y(_3305_));
 sky130_fd_sc_hd__nand3_1 _7350_ (.A(net82),
    .B(net99),
    .C(net100),
    .Y(_3306_));
 sky130_fd_sc_hd__or3b_1 _7351_ (.A(_3306_),
    .B(net405),
    .C_N(net393),
    .X(_3307_));
 sky130_fd_sc_hd__or2_1 _7352_ (.A(net397),
    .B(net411),
    .X(_3308_));
 sky130_fd_sc_hd__mux2_1 _7353_ (.A0(net447),
    .A1(\mul_wb.l[0] ),
    .S(net412),
    .X(_3309_));
 sky130_fd_sc_hd__and2_1 _7354_ (.A(net278),
    .B(net448),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _7355_ (.A0(net469),
    .A1(net485),
    .S(net412),
    .X(_3310_));
 sky130_fd_sc_hd__and2_1 _7356_ (.A(net278),
    .B(net486),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _7357_ (.A0(net481),
    .A1(net498),
    .S(net412),
    .X(_3311_));
 sky130_fd_sc_hd__and2_1 _7358_ (.A(net278),
    .B(net499),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _7359_ (.A0(net501),
    .A1(net512),
    .S(net412),
    .X(_3312_));
 sky130_fd_sc_hd__and2_1 _7360_ (.A(net278),
    .B(net513),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _7361_ (.A0(net474),
    .A1(\mul_wb.l[4] ),
    .S(net412),
    .X(_3313_));
 sky130_fd_sc_hd__and2_1 _7362_ (.A(net279),
    .B(net475),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _7363_ (.A0(net466),
    .A1(net478),
    .S(net412),
    .X(_3314_));
 sky130_fd_sc_hd__and2_1 _7364_ (.A(net279),
    .B(net479),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _7365_ (.A0(net463),
    .A1(net476),
    .S(net412),
    .X(_3315_));
 sky130_fd_sc_hd__and2_1 _7366_ (.A(net278),
    .B(net477),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _7367_ (.A0(net433),
    .A1(net437),
    .S(net412),
    .X(_3316_));
 sky130_fd_sc_hd__and2_1 _7368_ (.A(net279),
    .B(net438),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _7369_ (.A0(net415),
    .A1(net418),
    .S(net412),
    .X(_3317_));
 sky130_fd_sc_hd__and2_1 _7370_ (.A(net280),
    .B(net419),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _7371_ (.A0(net515),
    .A1(net522),
    .S(net412),
    .X(_3318_));
 sky130_fd_sc_hd__and2_1 _7372_ (.A(net279),
    .B(_3318_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _7373_ (.A0(net421),
    .A1(net424),
    .S(net412),
    .X(_3319_));
 sky130_fd_sc_hd__and2_1 _7374_ (.A(net280),
    .B(net425),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _7375_ (.A0(net401),
    .A1(\mul_wb.l[11] ),
    .S(net412),
    .X(_3320_));
 sky130_fd_sc_hd__and2_1 _7376_ (.A(net280),
    .B(net413),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _7377_ (.A0(net452),
    .A1(\mul_wb.l[12] ),
    .S(net412),
    .X(_3321_));
 sky130_fd_sc_hd__and2_1 _7378_ (.A(net280),
    .B(net453),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _7379_ (.A0(net488),
    .A1(net492),
    .S(net412),
    .X(_3322_));
 sky130_fd_sc_hd__and2_1 _7380_ (.A(net280),
    .B(net493),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _7381_ (.A0(net506),
    .A1(net510),
    .S(net412),
    .X(_3323_));
 sky130_fd_sc_hd__and2_1 _7382_ (.A(net280),
    .B(net511),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _7383_ (.A0(net440),
    .A1(\mul_wb.l[15] ),
    .S(net412),
    .X(_3324_));
 sky130_fd_sc_hd__and2_1 _7384_ (.A(_0000_),
    .B(net441),
    .X(_0176_));
 sky130_fd_sc_hd__nand2b_1 _7385_ (.A_N(net396),
    .B(net429),
    .Y(_3325_));
 sky130_fd_sc_hd__nand2_1 _7386_ (.A(net405),
    .B(net393),
    .Y(_3326_));
 sky130_fd_sc_hd__or3_1 _7387_ (.A(_3306_),
    .B(net430),
    .C(net406),
    .X(_3327_));
 sky130_fd_sc_hd__mux2_1 _7388_ (.A0(net447),
    .A1(net454),
    .S(net407),
    .X(_3328_));
 sky130_fd_sc_hd__and2_1 _7389_ (.A(net279),
    .B(net455),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _7390_ (.A0(net469),
    .A1(net471),
    .S(net407),
    .X(_3329_));
 sky130_fd_sc_hd__and2_1 _7391_ (.A(net278),
    .B(net472),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _7392_ (.A0(net481),
    .A1(\mul_wb.b[2] ),
    .S(net407),
    .X(_3330_));
 sky130_fd_sc_hd__and2_1 _7393_ (.A(net278),
    .B(net482),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _7394_ (.A0(net501),
    .A1(\mul_wb.b[3] ),
    .S(net407),
    .X(_3331_));
 sky130_fd_sc_hd__and2_1 _7395_ (.A(net279),
    .B(net502),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _7396_ (.A0(net474),
    .A1(net494),
    .S(net407),
    .X(_3332_));
 sky130_fd_sc_hd__and2_1 _7397_ (.A(net279),
    .B(net495),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _7398_ (.A0(net466),
    .A1(\mul_wb.b[5] ),
    .S(net407),
    .X(_3333_));
 sky130_fd_sc_hd__and2_1 _7399_ (.A(net279),
    .B(net467),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _7400_ (.A0(net463),
    .A1(net496),
    .S(net407),
    .X(_3334_));
 sky130_fd_sc_hd__and2_1 _7401_ (.A(net279),
    .B(net497),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _7402_ (.A0(net433),
    .A1(net449),
    .S(net407),
    .X(_3335_));
 sky130_fd_sc_hd__and2_1 _7403_ (.A(net279),
    .B(net450),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _7404_ (.A0(net415),
    .A1(\mul_wb.b[8] ),
    .S(net407),
    .X(_3336_));
 sky130_fd_sc_hd__and2_1 _7405_ (.A(net280),
    .B(net416),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _7406_ (.A0(net515),
    .A1(net521),
    .S(net407),
    .X(_3337_));
 sky130_fd_sc_hd__and2_1 _7407_ (.A(net280),
    .B(_3337_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _7408_ (.A0(net421),
    .A1(\mul_wb.b[10] ),
    .S(net407),
    .X(_3338_));
 sky130_fd_sc_hd__and2_1 _7409_ (.A(net280),
    .B(net422),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _7410_ (.A0(net401),
    .A1(\mul_wb.b[11] ),
    .S(net407),
    .X(_3339_));
 sky130_fd_sc_hd__and2_1 _7411_ (.A(net280),
    .B(net408),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _7412_ (.A0(net452),
    .A1(net460),
    .S(net407),
    .X(_3340_));
 sky130_fd_sc_hd__and2_1 _7413_ (.A(net280),
    .B(net461),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _7414_ (.A0(net488),
    .A1(\mul_wb.b[13] ),
    .S(net407),
    .X(_3341_));
 sky130_fd_sc_hd__and2_1 _7415_ (.A(_0000_),
    .B(net489),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _7416_ (.A0(net506),
    .A1(\mul_wb.b[14] ),
    .S(net407),
    .X(_3342_));
 sky130_fd_sc_hd__and2_1 _7417_ (.A(_0000_),
    .B(net507),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _7418_ (.A0(net440),
    .A1(net444),
    .S(net407),
    .X(_3343_));
 sky130_fd_sc_hd__and2_1 _7419_ (.A(net280),
    .B(net445),
    .X(_0192_));
 sky130_fd_sc_hd__or2_4 _7420_ (.A(net411),
    .B(net430),
    .X(_3344_));
 sky130_fd_sc_hd__mux2_1 _7421_ (.A0(net447),
    .A1(net458),
    .S(_3344_),
    .X(_3345_));
 sky130_fd_sc_hd__and2_1 _7422_ (.A(net279),
    .B(net459),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _7423_ (.A0(net469),
    .A1(\mul_wb.a[1] ),
    .S(_3344_),
    .X(_3346_));
 sky130_fd_sc_hd__and2_1 _7424_ (.A(net278),
    .B(net470),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _7425_ (.A0(net481),
    .A1(net503),
    .S(_3344_),
    .X(_3347_));
 sky130_fd_sc_hd__and2_1 _7426_ (.A(net278),
    .B(net504),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _7427_ (.A0(net501),
    .A1(net508),
    .S(_3344_),
    .X(_3348_));
 sky130_fd_sc_hd__and2_1 _7428_ (.A(net278),
    .B(net509),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _7429_ (.A0(net474),
    .A1(net490),
    .S(_3344_),
    .X(_3349_));
 sky130_fd_sc_hd__and2_1 _7430_ (.A(net278),
    .B(net491),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _7431_ (.A0(net466),
    .A1(net483),
    .S(_3344_),
    .X(_3350_));
 sky130_fd_sc_hd__and2_1 _7432_ (.A(net278),
    .B(net484),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _7433_ (.A0(net463),
    .A1(\mul_wb.a[6] ),
    .S(_3344_),
    .X(_3351_));
 sky130_fd_sc_hd__and2_1 _7434_ (.A(net278),
    .B(net464),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _7435_ (.A0(net433),
    .A1(\mul_wb.a[7] ),
    .S(_3344_),
    .X(_3352_));
 sky130_fd_sc_hd__and2_1 _7436_ (.A(net278),
    .B(net434),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _7437_ (.A0(net415),
    .A1(net435),
    .S(_3344_),
    .X(_3353_));
 sky130_fd_sc_hd__and2_1 _7438_ (.A(net279),
    .B(net436),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _7439_ (.A0(net515),
    .A1(\mul_wb.a[9] ),
    .S(_3344_),
    .X(_3354_));
 sky130_fd_sc_hd__and2_1 _7440_ (.A(net279),
    .B(net516),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _7441_ (.A0(net421),
    .A1(\mul_wb.a[10] ),
    .S(_3344_),
    .X(_3355_));
 sky130_fd_sc_hd__and2_1 _7442_ (.A(net280),
    .B(net431),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _7443_ (.A0(net401),
    .A1(\mul_wb.a[11] ),
    .S(_3344_),
    .X(_3356_));
 sky130_fd_sc_hd__and2_1 _7444_ (.A(net280),
    .B(net402),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _7445_ (.A0(net452),
    .A1(net456),
    .S(_3344_),
    .X(_3357_));
 sky130_fd_sc_hd__and2_1 _7446_ (.A(net280),
    .B(net457),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _7447_ (.A0(net488),
    .A1(net517),
    .S(_3344_),
    .X(_3358_));
 sky130_fd_sc_hd__and2_1 _7448_ (.A(_0000_),
    .B(net518),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _7449_ (.A0(net506),
    .A1(net519),
    .S(_3344_),
    .X(_3359_));
 sky130_fd_sc_hd__and2_1 _7450_ (.A(_0000_),
    .B(net520),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _7451_ (.A0(net440),
    .A1(net442),
    .S(_3344_),
    .X(_3360_));
 sky130_fd_sc_hd__and2_1 _7452_ (.A(net280),
    .B(net443),
    .X(_0208_));
 sky130_fd_sc_hd__nand3b_4 _7453_ (.A_N(net100),
    .B(net99),
    .C(net82),
    .Y(_3361_));
 sky130_fd_sc_hd__nor3_2 _7454_ (.A(net397),
    .B(net406),
    .C(net277),
    .Y(_3362_));
 sky130_fd_sc_hd__a22o_1 _7455_ (.A1(net134),
    .A2(net277),
    .B1(net230),
    .B2(net543),
    .X(_0209_));
 sky130_fd_sc_hd__a22o_1 _7456_ (.A1(net145),
    .A2(net277),
    .B1(net230),
    .B2(net545),
    .X(_0210_));
 sky130_fd_sc_hd__a22o_1 _7457_ (.A1(net156),
    .A2(net277),
    .B1(net230),
    .B2(net541),
    .X(_0211_));
 sky130_fd_sc_hd__a22o_1 _7458_ (.A1(net159),
    .A2(net277),
    .B1(net230),
    .B2(net531),
    .X(_0212_));
 sky130_fd_sc_hd__a22o_1 _7459_ (.A1(net160),
    .A2(net277),
    .B1(net230),
    .B2(net535),
    .X(_0213_));
 sky130_fd_sc_hd__a22o_1 _7460_ (.A1(net161),
    .A2(net277),
    .B1(net230),
    .B2(net533),
    .X(_0214_));
 sky130_fd_sc_hd__a22o_1 _7461_ (.A1(net162),
    .A2(net277),
    .B1(net230),
    .B2(net529),
    .X(_0215_));
 sky130_fd_sc_hd__a22o_1 _7462_ (.A1(net163),
    .A2(net277),
    .B1(net230),
    .B2(net547),
    .X(_0216_));
 sky130_fd_sc_hd__a22o_1 _7463_ (.A1(net164),
    .A2(net277),
    .B1(net230),
    .B2(net537),
    .X(_0217_));
 sky130_fd_sc_hd__a22o_1 _7464_ (.A1(net165),
    .A2(net277),
    .B1(net230),
    .B2(net525),
    .X(_0218_));
 sky130_fd_sc_hd__a22o_1 _7465_ (.A1(net135),
    .A2(net277),
    .B1(net230),
    .B2(net523),
    .X(_0219_));
 sky130_fd_sc_hd__a22o_1 _7466_ (.A1(net136),
    .A2(net277),
    .B1(net230),
    .B2(net539),
    .X(_0220_));
 sky130_fd_sc_hd__a22o_1 _7467_ (.A1(net137),
    .A2(net277),
    .B1(net230),
    .B2(net527),
    .X(_0221_));
 sky130_fd_sc_hd__a22o_1 _7468_ (.A1(net138),
    .A2(net276),
    .B1(net229),
    .B2(net617),
    .X(_0222_));
 sky130_fd_sc_hd__a22o_1 _7469_ (.A1(net139),
    .A2(net276),
    .B1(net229),
    .B2(net619),
    .X(_0223_));
 sky130_fd_sc_hd__a22o_1 _7470_ (.A1(net140),
    .A2(net276),
    .B1(net229),
    .B2(net621),
    .X(_0224_));
 sky130_fd_sc_hd__a22o_1 _7471_ (.A1(net141),
    .A2(net276),
    .B1(net229),
    .B2(net623),
    .X(_0225_));
 sky130_fd_sc_hd__a22o_1 _7472_ (.A1(net142),
    .A2(net276),
    .B1(net229),
    .B2(net629),
    .X(_0226_));
 sky130_fd_sc_hd__a22o_1 _7473_ (.A1(net143),
    .A2(net276),
    .B1(net229),
    .B2(net625),
    .X(_0227_));
 sky130_fd_sc_hd__a22o_1 _7474_ (.A1(net144),
    .A2(net276),
    .B1(net229),
    .B2(net627),
    .X(_0228_));
 sky130_fd_sc_hd__a22o_1 _7475_ (.A1(net146),
    .A2(net276),
    .B1(net229),
    .B2(net641),
    .X(_0229_));
 sky130_fd_sc_hd__a22o_1 _7476_ (.A1(net147),
    .A2(net276),
    .B1(net229),
    .B2(net631),
    .X(_0230_));
 sky130_fd_sc_hd__a22o_1 _7477_ (.A1(net148),
    .A2(net276),
    .B1(net229),
    .B2(net635),
    .X(_0231_));
 sky130_fd_sc_hd__a22o_1 _7478_ (.A1(net149),
    .A2(net276),
    .B1(net229),
    .B2(net637),
    .X(_0232_));
 sky130_fd_sc_hd__a22o_1 _7479_ (.A1(net150),
    .A2(net276),
    .B1(net229),
    .B2(net633),
    .X(_0233_));
 sky130_fd_sc_hd__a22o_1 _7480_ (.A1(net151),
    .A2(net276),
    .B1(net229),
    .B2(net645),
    .X(_0234_));
 sky130_fd_sc_hd__a22o_1 _7481_ (.A1(net152),
    .A2(net276),
    .B1(net229),
    .B2(net639),
    .X(_0235_));
 sky130_fd_sc_hd__a22o_1 _7482_ (.A1(net153),
    .A2(net276),
    .B1(net229),
    .B2(net647),
    .X(_0236_));
 sky130_fd_sc_hd__a22o_1 _7483_ (.A1(net154),
    .A2(net276),
    .B1(net229),
    .B2(net643),
    .X(_0237_));
 sky130_fd_sc_hd__a22o_1 _7484_ (.A1(net155),
    .A2(net277),
    .B1(net230),
    .B2(net615),
    .X(_0238_));
 sky130_fd_sc_hd__a22o_1 _7485_ (.A1(net157),
    .A2(_3361_),
    .B1(net230),
    .B2(net613),
    .X(_0239_));
 sky130_fd_sc_hd__a22o_1 _7486_ (.A1(net158),
    .A2(_3361_),
    .B1(net398),
    .B2(net991),
    .X(_0240_));
 sky130_fd_sc_hd__inv_2 _7487_ (.A(net281),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _7488_ (.A(net281),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _7489_ (.A(net281),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _7490_ (.A(net281),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _7491_ (.A(net281),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _7492_ (.A(net281),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _7493_ (.A(net281),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _7494_ (.A(net281),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _7495_ (.A(net281),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _7496_ (.A(net281),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _7497_ (.A(net281),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _7498_ (.A(net281),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _7499_ (.A(net283),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _7500_ (.A(net283),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _7501_ (.A(net285),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _7502_ (.A(net285),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _7503_ (.A(net285),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _7504_ (.A(net285),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _7505_ (.A(net285),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _7506_ (.A(net285),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _7507_ (.A(net285),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _7508_ (.A(net285),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _7509_ (.A(net285),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _7510_ (.A(net285),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _7511_ (.A(net286),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _7512_ (.A(net286),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _7513_ (.A(net287),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _7514_ (.A(net286),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _7515_ (.A(net286),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _7516_ (.A(net286),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _7517_ (.A(net286),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _7518_ (.A(net281),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _7519_ (.A(net282),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _7520_ (.A(net282),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _7521_ (.A(net282),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _7522_ (.A(net281),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _7523_ (.A(net282),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _7524_ (.A(net281),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _7525_ (.A(net282),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _7526_ (.A(net283),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _7527_ (.A(net284),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _7528_ (.A(net283),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _7529_ (.A(net283),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _7530_ (.A(net285),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _7531_ (.A(net286),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _7532_ (.A(net286),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _7533_ (.A(net285),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _7534_ (.A(net282),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _7535_ (.A(net282),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _7536_ (.A(net282),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _7537_ (.A(net283),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _7538_ (.A(net282),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _7539_ (.A(net283),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _7540_ (.A(net283),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _7541_ (.A(net283),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _7542_ (.A(net283),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _7543_ (.A(net283),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _7544_ (.A(net283),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _7545_ (.A(net283),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _7546_ (.A(net284),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _7547_ (.A(net285),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _7548_ (.A(net286),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _7549_ (.A(net285),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _7550_ (.A(net282),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _7551_ (.A(net282),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _7552_ (.A(net282),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _7553_ (.A(net282),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _7554_ (.A(net284),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _7555_ (.A(net284),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _7556_ (.A(net282),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _7557_ (.A(net282),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _7558_ (.A(net283),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _7559_ (.A(net284),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _7560_ (.A(net283),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _7561_ (.A(net283),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _7562_ (.A(net285),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _7563_ (.A(net284),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _7564_ (.A(net286),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _7565_ (.A(net285),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _7566_ (.A(net292),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _7567_ (.A(net292),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _7568_ (.A(net292),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _7569_ (.A(net292),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _7570_ (.A(net292),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _7571_ (.A(net292),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _7572_ (.A(net292),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _7573_ (.A(net292),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _7574_ (.A(net292),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _7575_ (.A(net290),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _7576_ (.A(net290),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _7577_ (.A(net290),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _7578_ (.A(net290),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _7579_ (.A(net290),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _7580_ (.A(net290),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _7581_ (.A(net290),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _7582_ (.A(net290),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _7583_ (.A(net290),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _7584_ (.A(net290),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _7585_ (.A(net290),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _7586_ (.A(net290),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _7587_ (.A(net290),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _7588_ (.A(net290),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _7589_ (.A(net290),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _7590_ (.A(net290),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _7591_ (.A(net291),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _7592_ (.A(net291),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _7593_ (.A(net291),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _7594_ (.A(net291),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _7595_ (.A(net291),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _7596_ (.A(net291),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _7597_ (.A(net291),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _7598_ (.A(net289),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _7599_ (.A(net289),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _7600_ (.A(net289),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _7601_ (.A(net289),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _7602_ (.A(net289),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _7603_ (.A(net289),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _7604_ (.A(net289),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _7605_ (.A(net289),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _7606_ (.A(net289),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _7607_ (.A(net292),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _7608_ (.A(net292),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _7609_ (.A(net292),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _7610_ (.A(net292),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _7611_ (.A(net292),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _7612_ (.A(net292),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _7613_ (.A(net292),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _7614_ (.A(net287),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _7615_ (.A(net287),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _7616_ (.A(net287),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _7617_ (.A(net288),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _7618_ (.A(net288),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _7619_ (.A(net288),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _7620_ (.A(net288),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _7621_ (.A(net289),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _7622_ (.A(net289),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _7623_ (.A(net289),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _7624_ (.A(net289),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _7625_ (.A(net289),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _7626_ (.A(net289),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _7627_ (.A(net289),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _7628_ (.A(net293),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _7629_ (.A(net293),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _7630_ (.A(net287),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _7631_ (.A(net287),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _7632_ (.A(net287),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _7633_ (.A(net287),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _7634_ (.A(net287),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _7635_ (.A(net287),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_2 _7636_ (.A(net287),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _7637_ (.A(net287),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _7638_ (.A(net287),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _7639_ (.A(net287),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _7640_ (.A(net287),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _7641_ (.A(net287),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _7642_ (.A(net288),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_2 _7643_ (.A(net288),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_2 _7644_ (.A(net288),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _7645_ (.A(net288),
    .Y(_0159_));
 sky130_fd_sc_hd__dfxtp_1 _7646_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net394),
    .Q(net133));
 sky130_fd_sc_hd__dfxtp_1 _7647_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0161_),
    .Q(\mul_wb.l[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7648_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0162_),
    .Q(\mul_wb.l[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7649_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0163_),
    .Q(\mul_wb.l[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7650_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0164_),
    .Q(\mul_wb.l[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7651_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0165_),
    .Q(\mul_wb.l[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7652_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0166_),
    .Q(\mul_wb.l[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7653_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0167_),
    .Q(\mul_wb.l[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7654_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0168_),
    .Q(\mul_wb.l[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7655_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0169_),
    .Q(\mul_wb.l[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7656_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0170_),
    .Q(\mul_wb.l[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7657_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0171_),
    .Q(\mul_wb.l[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7658_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0172_),
    .Q(\mul_wb.l[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7659_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0173_),
    .Q(\mul_wb.l[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7660_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0174_),
    .Q(\mul_wb.l[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7661_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0175_),
    .Q(\mul_wb.l[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7662_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0176_),
    .Q(\mul_wb.l[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7663_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0177_),
    .Q(\mul_wb.b[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7664_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0178_),
    .Q(\mul_wb.b[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7665_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0179_),
    .Q(\mul_wb.b[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7666_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0180_),
    .Q(\mul_wb.b[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7667_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0181_),
    .Q(\mul_wb.b[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7668_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0182_),
    .Q(\mul_wb.b[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7669_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0183_),
    .Q(\mul_wb.b[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7670_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0184_),
    .Q(\mul_wb.b[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7671_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net417),
    .Q(\mul_wb.b[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7672_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0186_),
    .Q(\mul_wb.b[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7673_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net423),
    .Q(\mul_wb.b[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7674_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net409),
    .Q(\mul_wb.b[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7675_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0189_),
    .Q(\mul_wb.b[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7676_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0190_),
    .Q(\mul_wb.b[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7677_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0191_),
    .Q(\mul_wb.b[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7678_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0192_),
    .Q(\mul_wb.b[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7679_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0193_),
    .Q(\mul_wb.a[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7680_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0194_),
    .Q(\mul_wb.a[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7681_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0195_),
    .Q(\mul_wb.a[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7682_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0196_),
    .Q(\mul_wb.a[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7683_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0197_),
    .Q(\mul_wb.a[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7684_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0198_),
    .Q(\mul_wb.a[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7685_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0199_),
    .Q(\mul_wb.a[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7686_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0200_),
    .Q(\mul_wb.a[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7687_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0201_),
    .Q(\mul_wb.a[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7688_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0202_),
    .Q(\mul_wb.a[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7689_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0203_),
    .Q(\mul_wb.a[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7690_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net403),
    .Q(\mul_wb.a[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7691_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0205_),
    .Q(\mul_wb.a[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7692_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0206_),
    .Q(\mul_wb.a[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7693_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0207_),
    .Q(\mul_wb.a[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7694_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0208_),
    .Q(\mul_wb.a[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7695_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net544),
    .Q(net134));
 sky130_fd_sc_hd__dfxtp_1 _7696_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net546),
    .Q(net145));
 sky130_fd_sc_hd__dfxtp_1 _7697_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net542),
    .Q(net156));
 sky130_fd_sc_hd__dfxtp_1 _7698_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net532),
    .Q(net159));
 sky130_fd_sc_hd__dfxtp_1 _7699_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net536),
    .Q(net160));
 sky130_fd_sc_hd__dfxtp_1 _7700_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net534),
    .Q(net161));
 sky130_fd_sc_hd__dfxtp_1 _7701_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net530),
    .Q(net162));
 sky130_fd_sc_hd__dfxtp_1 _7702_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net548),
    .Q(net163));
 sky130_fd_sc_hd__dfxtp_1 _7703_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net538),
    .Q(net164));
 sky130_fd_sc_hd__dfxtp_1 _7704_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net526),
    .Q(net165));
 sky130_fd_sc_hd__dfxtp_1 _7705_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net524),
    .Q(net135));
 sky130_fd_sc_hd__dfxtp_1 _7706_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net540),
    .Q(net136));
 sky130_fd_sc_hd__dfxtp_1 _7707_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net528),
    .Q(net137));
 sky130_fd_sc_hd__dfxtp_1 _7708_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net618),
    .Q(net138));
 sky130_fd_sc_hd__dfxtp_1 _7709_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net620),
    .Q(net139));
 sky130_fd_sc_hd__dfxtp_1 _7710_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net622),
    .Q(net140));
 sky130_fd_sc_hd__dfxtp_1 _7711_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net624),
    .Q(net141));
 sky130_fd_sc_hd__dfxtp_1 _7712_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net630),
    .Q(net142));
 sky130_fd_sc_hd__dfxtp_1 _7713_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net626),
    .Q(net143));
 sky130_fd_sc_hd__dfxtp_1 _7714_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net628),
    .Q(net144));
 sky130_fd_sc_hd__dfxtp_1 _7715_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net642),
    .Q(net146));
 sky130_fd_sc_hd__dfxtp_1 _7716_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net632),
    .Q(net147));
 sky130_fd_sc_hd__dfxtp_1 _7717_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net636),
    .Q(net148));
 sky130_fd_sc_hd__dfxtp_1 _7718_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net638),
    .Q(net149));
 sky130_fd_sc_hd__dfxtp_1 _7719_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net634),
    .Q(net150));
 sky130_fd_sc_hd__dfxtp_1 _7720_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net646),
    .Q(net151));
 sky130_fd_sc_hd__dfxtp_1 _7721_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net640),
    .Q(net152));
 sky130_fd_sc_hd__dfxtp_1 _7722_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net648),
    .Q(net153));
 sky130_fd_sc_hd__dfxtp_1 _7723_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net644),
    .Q(net154));
 sky130_fd_sc_hd__dfxtp_1 _7724_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net616),
    .Q(net155));
 sky130_fd_sc_hd__dfxtp_1 _7725_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net614),
    .Q(net157));
 sky130_fd_sc_hd__dfxtp_1 _7726_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net399),
    .Q(net158));
 sky130_fd_sc_hd__dfrtp_1 _7727_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(\mul_wb.P_[0] ),
    .RESET_B(net278),
    .Q(\mul_wb.p[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7728_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(\mul_wb.reg_p[1] ),
    .RESET_B(_0001_),
    .Q(\mul_wb.p[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7729_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(\mul_wb.reg_p[2] ),
    .RESET_B(_0002_),
    .Q(\mul_wb.p[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7730_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\mul_wb.reg_p[3] ),
    .RESET_B(_0003_),
    .Q(\mul_wb.p[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7731_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(\mul_wb.reg_p[4] ),
    .RESET_B(_0004_),
    .Q(\mul_wb.p[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7732_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\mul_wb.reg_p[5] ),
    .RESET_B(_0005_),
    .Q(\mul_wb.p[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7733_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\mul_wb.reg_p[6] ),
    .RESET_B(_0006_),
    .Q(\mul_wb.p[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7734_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\mul_wb.reg_p[7] ),
    .RESET_B(_0007_),
    .Q(\mul_wb.p[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7735_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\mul_wb.reg_p[8] ),
    .RESET_B(_0008_),
    .Q(\mul_wb.p[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7736_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\mul_wb.reg_p[9] ),
    .RESET_B(_0009_),
    .Q(\mul_wb.p[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7737_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\mul_wb.reg_p[10] ),
    .RESET_B(_0010_),
    .Q(\mul_wb.p[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7738_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\mul_wb.reg_p[11] ),
    .RESET_B(_0011_),
    .Q(\mul_wb.p[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7739_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(\mul_wb.reg_p[12] ),
    .RESET_B(_0012_),
    .Q(\mul_wb.p[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7740_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(\mul_wb.reg_p[13] ),
    .RESET_B(_0013_),
    .Q(\mul_wb.p[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7741_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(\mul_wb.reg_p[14] ),
    .RESET_B(_0014_),
    .Q(\mul_wb.p[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7742_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(\mul_wb.reg_p[15] ),
    .RESET_B(_0015_),
    .Q(\mul_wb.p[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7743_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(\mul_wb.reg_p[16] ),
    .RESET_B(_0016_),
    .Q(\mul_wb.p[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7744_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(\mul_wb.reg_p[17] ),
    .RESET_B(_0017_),
    .Q(\mul_wb.p[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7745_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(\mul_wb.reg_p[18] ),
    .RESET_B(_0018_),
    .Q(\mul_wb.p[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7746_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(\mul_wb.reg_p[19] ),
    .RESET_B(_0019_),
    .Q(\mul_wb.p[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7747_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(\mul_wb.reg_p[20] ),
    .RESET_B(_0020_),
    .Q(\mul_wb.p[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7748_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(\mul_wb.reg_p[21] ),
    .RESET_B(_0021_),
    .Q(\mul_wb.p[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7749_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(\mul_wb.reg_p[22] ),
    .RESET_B(_0022_),
    .Q(\mul_wb.p[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7750_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(\mul_wb.reg_p[23] ),
    .RESET_B(_0023_),
    .Q(\mul_wb.p[23] ));
 sky130_fd_sc_hd__dfrtp_1 _7751_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(\mul_wb.reg_p[24] ),
    .RESET_B(_0024_),
    .Q(\mul_wb.p[24] ));
 sky130_fd_sc_hd__dfrtp_1 _7752_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(\mul_wb.reg_p[25] ),
    .RESET_B(_0025_),
    .Q(\mul_wb.p[25] ));
 sky130_fd_sc_hd__dfrtp_1 _7753_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(\mul_wb.reg_p[26] ),
    .RESET_B(_0026_),
    .Q(\mul_wb.p[26] ));
 sky130_fd_sc_hd__dfrtp_1 _7754_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(\mul_wb.reg_p[27] ),
    .RESET_B(_0027_),
    .Q(\mul_wb.p[27] ));
 sky130_fd_sc_hd__dfrtp_1 _7755_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(\mul_wb.reg_p[28] ),
    .RESET_B(_0028_),
    .Q(\mul_wb.p[28] ));
 sky130_fd_sc_hd__dfrtp_1 _7756_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(\mul_wb.reg_p[29] ),
    .RESET_B(_0029_),
    .Q(\mul_wb.p[29] ));
 sky130_fd_sc_hd__dfrtp_1 _7757_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(\mul_wb.reg_p[30] ),
    .RESET_B(_0030_),
    .Q(\mul_wb.p[30] ));
 sky130_fd_sc_hd__dfrtp_1 _7758_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(\mul_wb.reg_p[31] ),
    .RESET_B(_0031_),
    .Q(\mul_wb.p[31] ));
 sky130_fd_sc_hd__dfrtp_2 _7759_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net672),
    .RESET_B(_0032_),
    .Q(\mul_wb.lob_4.L[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7760_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net485),
    .RESET_B(_0033_),
    .Q(\mul_wb.lob_4.L[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7761_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net498),
    .RESET_B(_0034_),
    .Q(\mul_wb.lob_4.L[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7762_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net512),
    .RESET_B(_0035_),
    .Q(\mul_wb.lob_4.L[3] ));
 sky130_fd_sc_hd__dfrtp_4 _7763_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net657),
    .RESET_B(_0036_),
    .Q(\mul_wb.lob_4.L[4] ));
 sky130_fd_sc_hd__dfrtp_4 _7764_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net478),
    .RESET_B(_0037_),
    .Q(\mul_wb.lob_4.L[5] ));
 sky130_fd_sc_hd__dfrtp_4 _7765_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net476),
    .RESET_B(_0038_),
    .Q(\mul_wb.lob_4.L[6] ));
 sky130_fd_sc_hd__dfrtp_4 _7766_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net437),
    .RESET_B(_0039_),
    .Q(\mul_wb.lob_4.L[7] ));
 sky130_fd_sc_hd__dfrtp_4 _7767_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net418),
    .RESET_B(_0040_),
    .Q(\mul_wb.lob_4.L[8] ));
 sky130_fd_sc_hd__dfrtp_4 _7768_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net522),
    .RESET_B(_0041_),
    .Q(\mul_wb.lob_4.L[9] ));
 sky130_fd_sc_hd__dfrtp_2 _7769_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net424),
    .RESET_B(_0042_),
    .Q(\mul_wb.lob_4.L[10] ));
 sky130_fd_sc_hd__dfrtp_2 _7770_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net691),
    .RESET_B(_0043_),
    .Q(\mul_wb.lob_4.L[11] ));
 sky130_fd_sc_hd__dfrtp_4 _7771_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net662),
    .RESET_B(_0044_),
    .Q(\mul_wb.lob_4.L[12] ));
 sky130_fd_sc_hd__dfrtp_4 _7772_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net492),
    .RESET_B(_0045_),
    .Q(\mul_wb.lob_4.L[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7773_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net510),
    .RESET_B(_0046_),
    .Q(\mul_wb.lob_4.L[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7774_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net692),
    .RESET_B(_0047_),
    .Q(\mul_wb.lob_4.L[15] ));
 sky130_fd_sc_hd__dfrtp_4 _7775_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net454),
    .RESET_B(_0048_),
    .Q(\mul_wb.lob_4.B[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7776_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net471),
    .RESET_B(_0049_),
    .Q(\mul_wb.reg_b0[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7777_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net687),
    .RESET_B(_0050_),
    .Q(\mul_wb.reg_b0[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7778_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net668),
    .RESET_B(_0051_),
    .Q(\mul_wb.reg_b0[3] ));
 sky130_fd_sc_hd__dfrtp_4 _7779_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net494),
    .RESET_B(_0052_),
    .Q(\mul_wb.reg_b0[4] ));
 sky130_fd_sc_hd__dfrtp_4 _7780_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net660),
    .RESET_B(_0053_),
    .Q(\mul_wb.reg_b0[5] ));
 sky130_fd_sc_hd__dfrtp_4 _7781_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net496),
    .RESET_B(_0054_),
    .Q(\mul_wb.reg_b0[6] ));
 sky130_fd_sc_hd__dfrtp_4 _7782_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net449),
    .RESET_B(_0055_),
    .Q(\mul_wb.reg_b0[7] ));
 sky130_fd_sc_hd__dfrtp_4 _7783_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net659),
    .RESET_B(_0056_),
    .Q(\mul_wb.reg_b0[8] ));
 sky130_fd_sc_hd__dfrtp_4 _7784_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net521),
    .RESET_B(_0057_),
    .Q(\mul_wb.reg_b0[9] ));
 sky130_fd_sc_hd__dfrtp_4 _7785_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net656),
    .RESET_B(_0058_),
    .Q(\mul_wb.reg_b0[10] ));
 sky130_fd_sc_hd__dfrtp_4 _7786_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net685),
    .RESET_B(_0059_),
    .Q(\mul_wb.reg_b0[11] ));
 sky130_fd_sc_hd__dfrtp_2 _7787_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net460),
    .RESET_B(_0060_),
    .Q(\mul_wb.reg_b0[12] ));
 sky130_fd_sc_hd__dfrtp_4 _7788_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net688),
    .RESET_B(_0061_),
    .Q(\mul_wb.reg_b0[13] ));
 sky130_fd_sc_hd__dfrtp_4 _7789_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net686),
    .RESET_B(_0062_),
    .Q(\mul_wb.reg_b0[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7790_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net444),
    .RESET_B(_0063_),
    .Q(\mul_wb.reg_b0[15] ));
 sky130_fd_sc_hd__dfrtp_4 _7791_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net458),
    .RESET_B(_0064_),
    .Q(\mul_wb.lob_4.A[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7792_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net666),
    .RESET_B(_0065_),
    .Q(\mul_wb.reg_a0[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7793_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net503),
    .RESET_B(_0066_),
    .Q(\mul_wb.reg_a0[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7794_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net508),
    .RESET_B(_0067_),
    .Q(\mul_wb.reg_a0[3] ));
 sky130_fd_sc_hd__dfrtp_4 _7795_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net490),
    .RESET_B(_0068_),
    .Q(\mul_wb.reg_a0[4] ));
 sky130_fd_sc_hd__dfrtp_2 _7796_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net483),
    .RESET_B(_0069_),
    .Q(\mul_wb.reg_a0[5] ));
 sky130_fd_sc_hd__dfrtp_4 _7797_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net670),
    .RESET_B(_0070_),
    .Q(\mul_wb.reg_a0[6] ));
 sky130_fd_sc_hd__dfrtp_4 _7798_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net678),
    .RESET_B(_0071_),
    .Q(\mul_wb.reg_a0[7] ));
 sky130_fd_sc_hd__dfrtp_4 _7799_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net435),
    .RESET_B(_0072_),
    .Q(\mul_wb.reg_a0[8] ));
 sky130_fd_sc_hd__dfrtp_4 _7800_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net665),
    .RESET_B(_0073_),
    .Q(\mul_wb.reg_a0[9] ));
 sky130_fd_sc_hd__dfrtp_4 _7801_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net694),
    .RESET_B(_0074_),
    .Q(\mul_wb.reg_a0[10] ));
 sky130_fd_sc_hd__dfrtp_2 _7802_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net696),
    .RESET_B(_0075_),
    .Q(\mul_wb.reg_a0[11] ));
 sky130_fd_sc_hd__dfrtp_4 _7803_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net456),
    .RESET_B(_0076_),
    .Q(\mul_wb.reg_a0[12] ));
 sky130_fd_sc_hd__dfrtp_4 _7804_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net517),
    .RESET_B(_0077_),
    .Q(\mul_wb.reg_a0[13] ));
 sky130_fd_sc_hd__dfrtp_4 _7805_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net519),
    .RESET_B(_0078_),
    .Q(\mul_wb.reg_a0[14] ));
 sky130_fd_sc_hd__dfrtp_2 _7806_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net442),
    .RESET_B(_0079_),
    .Q(\mul_wb.reg_a0[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7807_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(\mul_la.P_[0] ),
    .RESET_B(_0080_),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_1 _7808_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(\mul_la.reg_p[1] ),
    .RESET_B(_0081_),
    .Q(net112));
 sky130_fd_sc_hd__dfrtp_1 _7809_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(\mul_la.reg_p[2] ),
    .RESET_B(_0082_),
    .Q(net123));
 sky130_fd_sc_hd__dfrtp_1 _7810_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(\mul_la.reg_p[3] ),
    .RESET_B(_0083_),
    .Q(net126));
 sky130_fd_sc_hd__dfrtp_1 _7811_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(\mul_la.reg_p[4] ),
    .RESET_B(_0084_),
    .Q(net127));
 sky130_fd_sc_hd__dfrtp_1 _7812_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(\mul_la.reg_p[5] ),
    .RESET_B(_0085_),
    .Q(net128));
 sky130_fd_sc_hd__dfrtp_1 _7813_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(\mul_la.reg_p[6] ),
    .RESET_B(_0086_),
    .Q(net129));
 sky130_fd_sc_hd__dfrtp_1 _7814_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(\mul_la.reg_p[7] ),
    .RESET_B(_0087_),
    .Q(net130));
 sky130_fd_sc_hd__dfrtp_1 _7815_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\mul_la.reg_p[8] ),
    .RESET_B(_0088_),
    .Q(net131));
 sky130_fd_sc_hd__dfrtp_1 _7816_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\mul_la.reg_p[9] ),
    .RESET_B(_0089_),
    .Q(net132));
 sky130_fd_sc_hd__dfrtp_1 _7817_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\mul_la.reg_p[10] ),
    .RESET_B(_0090_),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_1 _7818_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\mul_la.reg_p[11] ),
    .RESET_B(_0091_),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_1 _7819_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\mul_la.reg_p[12] ),
    .RESET_B(_0092_),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_1 _7820_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\mul_la.reg_p[13] ),
    .RESET_B(_0093_),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_1 _7821_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\mul_la.reg_p[14] ),
    .RESET_B(_0094_),
    .Q(net106));
 sky130_fd_sc_hd__dfrtp_1 _7822_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\mul_la.reg_p[15] ),
    .RESET_B(_0095_),
    .Q(net107));
 sky130_fd_sc_hd__dfrtp_1 _7823_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\mul_la.reg_p[16] ),
    .RESET_B(_0096_),
    .Q(net108));
 sky130_fd_sc_hd__dfrtp_1 _7824_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\mul_la.reg_p[17] ),
    .RESET_B(_0097_),
    .Q(net109));
 sky130_fd_sc_hd__dfrtp_1 _7825_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\mul_la.reg_p[18] ),
    .RESET_B(_0098_),
    .Q(net110));
 sky130_fd_sc_hd__dfrtp_1 _7826_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\mul_la.reg_p[19] ),
    .RESET_B(_0099_),
    .Q(net111));
 sky130_fd_sc_hd__dfrtp_1 _7827_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\mul_la.reg_p[20] ),
    .RESET_B(_0100_),
    .Q(net113));
 sky130_fd_sc_hd__dfrtp_1 _7828_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\mul_la.reg_p[21] ),
    .RESET_B(_0101_),
    .Q(net114));
 sky130_fd_sc_hd__dfrtp_1 _7829_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\mul_la.reg_p[22] ),
    .RESET_B(_0102_),
    .Q(net115));
 sky130_fd_sc_hd__dfrtp_1 _7830_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\mul_la.reg_p[23] ),
    .RESET_B(_0103_),
    .Q(net116));
 sky130_fd_sc_hd__dfrtp_1 _7831_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\mul_la.reg_p[24] ),
    .RESET_B(_0104_),
    .Q(net117));
 sky130_fd_sc_hd__dfrtp_1 _7832_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\mul_la.reg_p[25] ),
    .RESET_B(_0105_),
    .Q(net118));
 sky130_fd_sc_hd__dfrtp_1 _7833_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\mul_la.reg_p[26] ),
    .RESET_B(_0106_),
    .Q(net119));
 sky130_fd_sc_hd__dfrtp_1 _7834_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\mul_la.reg_p[27] ),
    .RESET_B(_0107_),
    .Q(net120));
 sky130_fd_sc_hd__dfrtp_1 _7835_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\mul_la.reg_p[28] ),
    .RESET_B(_0108_),
    .Q(net121));
 sky130_fd_sc_hd__dfrtp_1 _7836_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\mul_la.reg_p[29] ),
    .RESET_B(_0109_),
    .Q(net122));
 sky130_fd_sc_hd__dfrtp_1 _7837_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net708),
    .RESET_B(_0110_),
    .Q(net124));
 sky130_fd_sc_hd__dfrtp_1 _7838_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(\mul_la.reg_p[31] ),
    .RESET_B(_0111_),
    .Q(net125));
 sky130_fd_sc_hd__dfrtp_2 _7839_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net813),
    .RESET_B(_0112_),
    .Q(\mul_la.lob_4.L[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7840_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net877),
    .RESET_B(_0113_),
    .Q(\mul_la.lob_4.L[1] ));
 sky130_fd_sc_hd__dfrtp_2 _7841_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net753),
    .RESET_B(_0114_),
    .Q(\mul_la.lob_4.L[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7842_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net713),
    .RESET_B(_0115_),
    .Q(\mul_la.lob_4.L[3] ));
 sky130_fd_sc_hd__dfrtp_4 _7843_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net745),
    .RESET_B(_0116_),
    .Q(\mul_la.lob_4.L[4] ));
 sky130_fd_sc_hd__dfrtp_4 _7844_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net729),
    .RESET_B(_0117_),
    .Q(\mul_la.lob_4.L[5] ));
 sky130_fd_sc_hd__dfrtp_4 _7845_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net721),
    .RESET_B(_0118_),
    .Q(\mul_la.lob_4.L[6] ));
 sky130_fd_sc_hd__dfrtp_4 _7846_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net737),
    .RESET_B(_0119_),
    .Q(\mul_la.lob_4.L[7] ));
 sky130_fd_sc_hd__dfrtp_4 _7847_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net761),
    .RESET_B(_0120_),
    .Q(\mul_la.lob_4.L[8] ));
 sky130_fd_sc_hd__dfrtp_2 _7848_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net717),
    .RESET_B(_0121_),
    .Q(\mul_la.lob_4.L[9] ));
 sky130_fd_sc_hd__dfrtp_4 _7849_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net789),
    .RESET_B(_0122_),
    .Q(\mul_la.lob_4.L[10] ));
 sky130_fd_sc_hd__dfrtp_4 _7850_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net733),
    .RESET_B(_0123_),
    .Q(\mul_la.lob_4.L[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7851_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net849),
    .RESET_B(_0124_),
    .Q(\mul_la.lob_4.L[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7852_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net841),
    .RESET_B(_0125_),
    .Q(\mul_la.lob_4.L[13] ));
 sky130_fd_sc_hd__dfrtp_2 _7853_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net749),
    .RESET_B(_0126_),
    .Q(\mul_la.lob_4.L[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7854_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net805),
    .RESET_B(_0127_),
    .Q(\mul_la.lob_4.L[15] ));
 sky130_fd_sc_hd__dfrtp_4 _7855_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net865),
    .RESET_B(_0128_),
    .Q(\mul_la.lob_4.B[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7856_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net793),
    .RESET_B(_0129_),
    .Q(\mul_la.reg_b0[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7857_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net769),
    .RESET_B(_0130_),
    .Q(\mul_la.reg_b0[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7858_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net817),
    .RESET_B(_0131_),
    .Q(\mul_la.reg_b0[3] ));
 sky130_fd_sc_hd__dfrtp_4 _7859_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net773),
    .RESET_B(_0132_),
    .Q(\mul_la.reg_b0[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7860_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net861),
    .RESET_B(_0133_),
    .Q(\mul_la.reg_b0[5] ));
 sky130_fd_sc_hd__dfrtp_4 _7861_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net845),
    .RESET_B(_0134_),
    .Q(\mul_la.reg_b0[6] ));
 sky130_fd_sc_hd__dfrtp_4 _7862_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net821),
    .RESET_B(_0135_),
    .Q(\mul_la.reg_b0[7] ));
 sky130_fd_sc_hd__dfrtp_4 _7863_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net825),
    .RESET_B(_0136_),
    .Q(\mul_la.reg_b0[8] ));
 sky130_fd_sc_hd__dfrtp_4 _7864_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net829),
    .RESET_B(_0137_),
    .Q(\mul_la.reg_b0[9] ));
 sky130_fd_sc_hd__dfrtp_4 _7865_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net809),
    .RESET_B(_0138_),
    .Q(\mul_la.reg_b0[10] ));
 sky130_fd_sc_hd__dfrtp_4 _7866_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net797),
    .RESET_B(_0139_),
    .Q(\mul_la.reg_b0[11] ));
 sky130_fd_sc_hd__dfrtp_4 _7867_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net857),
    .RESET_B(_0140_),
    .Q(\mul_la.reg_b0[12] ));
 sky130_fd_sc_hd__dfrtp_4 _7868_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net837),
    .RESET_B(_0141_),
    .Q(\mul_la.reg_b0[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7869_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net853),
    .RESET_B(_0142_),
    .Q(\mul_la.reg_b0[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7870_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net833),
    .RESET_B(_0143_),
    .Q(\mul_la.reg_b0[15] ));
 sky130_fd_sc_hd__dfrtp_4 _7871_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net897),
    .RESET_B(_0144_),
    .Q(\mul_la.lob_4.A[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7872_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net889),
    .RESET_B(_0145_),
    .Q(\mul_la.reg_a0[1] ));
 sky130_fd_sc_hd__dfrtp_2 _7873_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net901),
    .RESET_B(_0146_),
    .Q(\mul_la.reg_a0[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7874_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net893),
    .RESET_B(_0147_),
    .Q(\mul_la.reg_a0[3] ));
 sky130_fd_sc_hd__dfrtp_4 _7875_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net869),
    .RESET_B(_0148_),
    .Q(\mul_la.reg_a0[4] ));
 sky130_fd_sc_hd__dfrtp_4 _7876_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net885),
    .RESET_B(_0149_),
    .Q(\mul_la.reg_a0[5] ));
 sky130_fd_sc_hd__dfrtp_4 _7877_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net873),
    .RESET_B(_0150_),
    .Q(\mul_la.reg_a0[6] ));
 sky130_fd_sc_hd__dfrtp_4 _7878_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net881),
    .RESET_B(_0151_),
    .Q(\mul_la.reg_a0[7] ));
 sky130_fd_sc_hd__dfrtp_2 _7879_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net765),
    .RESET_B(_0152_),
    .Q(\mul_la.reg_a0[8] ));
 sky130_fd_sc_hd__dfrtp_4 _7880_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net757),
    .RESET_B(_0153_),
    .Q(\mul_la.reg_a0[9] ));
 sky130_fd_sc_hd__dfrtp_4 _7881_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net725),
    .RESET_B(_0154_),
    .Q(\mul_la.reg_a0[10] ));
 sky130_fd_sc_hd__dfrtp_2 _7882_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net801),
    .RESET_B(_0155_),
    .Q(\mul_la.reg_a0[11] ));
 sky130_fd_sc_hd__dfrtp_4 _7883_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net741),
    .RESET_B(_0156_),
    .Q(\mul_la.reg_a0[12] ));
 sky130_fd_sc_hd__dfrtp_4 _7884_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net777),
    .RESET_B(_0157_),
    .Q(\mul_la.reg_a0[13] ));
 sky130_fd_sc_hd__dfrtp_4 _7885_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net781),
    .RESET_B(_0158_),
    .Q(\mul_la.reg_a0[14] ));
 sky130_fd_sc_hd__dfrtp_4 _7886_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net785),
    .RESET_B(_0159_),
    .Q(\mul_la.reg_a0[15] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__buf_4 fanout167 (.A(_1775_),
    .X(net167));
 sky130_fd_sc_hd__buf_4 fanout168 (.A(_1979_),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_8 fanout169 (.A(_1934_),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_8 fanout170 (.A(net171),
    .X(net170));
 sky130_fd_sc_hd__buf_4 fanout172 (.A(_1828_),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_8 fanout173 (.A(_3657_),
    .X(net173));
 sky130_fd_sc_hd__buf_4 fanout174 (.A(_3587_),
    .X(net174));
 sky130_fd_sc_hd__buf_4 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_4 fanout176 (.A(_3562_),
    .X(net176));
 sky130_fd_sc_hd__buf_6 fanout177 (.A(_3475_),
    .X(net177));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(_2377_),
    .X(net178));
 sky130_fd_sc_hd__buf_6 fanout179 (.A(_2303_),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_8 fanout181 (.A(_2115_),
    .X(net181));
 sky130_fd_sc_hd__buf_4 fanout182 (.A(_2085_),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_2 fanout183 (.A(_2085_),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_8 fanout186 (.A(_1914_),
    .X(net186));
 sky130_fd_sc_hd__buf_4 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__buf_2 fanout188 (.A(_1663_),
    .X(net188));
 sky130_fd_sc_hd__buf_4 fanout189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_8 fanout190 (.A(_0503_),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_8 fanout191 (.A(_0442_),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_8 fanout192 (.A(_0399_),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_4 fanout193 (.A(_0399_),
    .X(net193));
 sky130_fd_sc_hd__buf_4 fanout194 (.A(_0391_),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_8 fanout195 (.A(_0346_),
    .X(net195));
 sky130_fd_sc_hd__buf_4 fanout196 (.A(_0332_),
    .X(net196));
 sky130_fd_sc_hd__buf_4 fanout197 (.A(_0332_),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_8 fanout198 (.A(_0286_),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_4 fanout199 (.A(_0286_),
    .X(net199));
 sky130_fd_sc_hd__buf_4 fanout200 (.A(_0272_),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_4 fanout201 (.A(_0272_),
    .X(net201));
 sky130_fd_sc_hd__buf_4 fanout202 (.A(_3783_),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_4 fanout203 (.A(_3783_),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_8 fanout204 (.A(_3773_),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_8 fanout206 (.A(_3722_),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_8 fanout207 (.A(_3697_),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_8 fanout208 (.A(_3683_),
    .X(net208));
 sky130_fd_sc_hd__buf_4 fanout209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_4 fanout210 (.A(_3641_),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_8 fanout213 (.A(_2234_),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_8 fanout214 (.A(_2175_),
    .X(net214));
 sky130_fd_sc_hd__buf_4 fanout216 (.A(_0753_),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_8 fanout217 (.A(_0715_),
    .X(net217));
 sky130_fd_sc_hd__buf_4 fanout218 (.A(_0637_),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_4 fanout219 (.A(_0637_),
    .X(net219));
 sky130_fd_sc_hd__buf_4 fanout220 (.A(_0607_),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_8 fanout221 (.A(_0598_),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_8 fanout222 (.A(_0535_),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_8 fanout223 (.A(_0472_),
    .X(net223));
 sky130_fd_sc_hd__buf_2 fanout224 (.A(_0472_),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_8 fanout225 (.A(_2524_),
    .X(net225));
 sky130_fd_sc_hd__buf_4 fanout227 (.A(_0667_),
    .X(net227));
 sky130_fd_sc_hd__buf_4 fanout229 (.A(net230),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_8 fanout230 (.A(net398),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_8 fanout232 (.A(_1693_),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_8 fanout233 (.A(_1692_),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_4 fanout235 (.A(_1599_),
    .X(net235));
 sky130_fd_sc_hd__buf_4 fanout236 (.A(_1577_),
    .X(net236));
 sky130_fd_sc_hd__buf_4 fanout237 (.A(_0816_),
    .X(net237));
 sky130_fd_sc_hd__buf_4 fanout243 (.A(_3493_),
    .X(net243));
 sky130_fd_sc_hd__buf_4 fanout244 (.A(_3484_),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_8 fanout246 (.A(_3401_),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_8 fanout248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_4 fanout249 (.A(_3395_),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_8 fanout250 (.A(_3390_),
    .X(net250));
 sky130_fd_sc_hd__buf_4 fanout251 (.A(net700),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_8 fanout252 (.A(net698),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_8 fanout253 (.A(\mul_la.reg_a0[15] ),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_8 fanout254 (.A(\mul_la.reg_b0[15] ),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_8 fanout255 (.A(net256),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_8 fanout256 (.A(\mul_la.lob_4.L[15] ),
    .X(net256));
 sky130_fd_sc_hd__buf_4 fanout257 (.A(\mul_la.lob_4.L[14] ),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_4 fanout258 (.A(\mul_la.lob_4.L[14] ),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_8 fanout259 (.A(\mul_la.lob_4.L[13] ),
    .X(net259));
 sky130_fd_sc_hd__buf_2 fanout260 (.A(\mul_la.lob_4.L[13] ),
    .X(net260));
 sky130_fd_sc_hd__buf_4 fanout261 (.A(\mul_la.lob_4.L[12] ),
    .X(net261));
 sky130_fd_sc_hd__buf_2 fanout262 (.A(\mul_la.lob_4.L[12] ),
    .X(net262));
 sky130_fd_sc_hd__buf_4 fanout263 (.A(\mul_la.lob_4.L[11] ),
    .X(net263));
 sky130_fd_sc_hd__buf_4 fanout264 (.A(\mul_la.lob_4.L[10] ),
    .X(net264));
 sky130_fd_sc_hd__buf_4 fanout265 (.A(\mul_la.lob_4.L[9] ),
    .X(net265));
 sky130_fd_sc_hd__buf_4 fanout266 (.A(\mul_wb.reg_a0[15] ),
    .X(net266));
 sky130_fd_sc_hd__buf_6 fanout267 (.A(net697),
    .X(net267));
 sky130_fd_sc_hd__buf_6 fanout268 (.A(\mul_wb.lob_4.L[15] ),
    .X(net268));
 sky130_fd_sc_hd__buf_8 fanout269 (.A(net701),
    .X(net269));
 sky130_fd_sc_hd__buf_4 fanout270 (.A(\mul_wb.lob_4.L[14] ),
    .X(net270));
 sky130_fd_sc_hd__buf_2 fanout271 (.A(\mul_wb.lob_4.L[14] ),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_8 fanout272 (.A(\mul_wb.lob_4.L[13] ),
    .X(net272));
 sky130_fd_sc_hd__buf_4 fanout273 (.A(\mul_wb.lob_4.L[12] ),
    .X(net273));
 sky130_fd_sc_hd__buf_4 fanout274 (.A(\mul_wb.lob_4.L[11] ),
    .X(net274));
 sky130_fd_sc_hd__buf_4 fanout275 (.A(\mul_wb.lob_4.L[10] ),
    .X(net275));
 sky130_fd_sc_hd__buf_4 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__buf_6 fanout277 (.A(_3361_),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_4 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_4 fanout279 (.A(_0000_),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_4 fanout280 (.A(_0000_),
    .X(net280));
 sky130_fd_sc_hd__buf_8 fanout281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__buf_8 fanout282 (.A(net284),
    .X(net282));
 sky130_fd_sc_hd__buf_8 fanout283 (.A(net284),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_8 fanout284 (.A(net293),
    .X(net284));
 sky130_fd_sc_hd__buf_8 fanout285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_8 fanout286 (.A(net293),
    .X(net286));
 sky130_fd_sc_hd__buf_8 fanout287 (.A(net293),
    .X(net287));
 sky130_fd_sc_hd__buf_4 fanout288 (.A(net293),
    .X(net288));
 sky130_fd_sc_hd__buf_8 fanout289 (.A(net293),
    .X(net289));
 sky130_fd_sc_hd__buf_8 fanout290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__buf_4 fanout291 (.A(net293),
    .X(net291));
 sky130_fd_sc_hd__buf_6 fanout292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__buf_8 fanout293 (.A(net49),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net714),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net736),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_0160_),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(wbs_adr_i[3]),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(net75),
    .X(net396));
 sky130_fd_sc_hd__buf_1 hold103 (.A(_3305_),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_2 hold104 (.A(_3362_),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_0240_),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(wbs_dat_i[11]),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(net85),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_3356_),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0204_),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net798),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(wbs_adr_i[2]),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(net72),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_3326_),
    .X(net406));
 sky130_fd_sc_hd__buf_6 hold113 (.A(_3327_),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_3339_),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_0188_),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(wbs_adr_i[0]),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_3307_),
    .X(net411));
 sky130_fd_sc_hd__buf_6 hold118 (.A(_3308_),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_3320_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net800),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(wbs_dat_i[8]),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(net97),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_3336_),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_0185_),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(net684),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_3317_),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(wbs_dat_i[10]),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(net84),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_3338_),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_0187_),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net770),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(net681),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_3319_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(wbs_adr_i[26]),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(net68),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_3296_),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_2 hold135 (.A(net968),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_3325_),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_3355_),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(wbs_dat_i[7]),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(net96),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net772),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_3352_),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(net651),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_3353_),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(net679),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_3316_),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(wbs_dat_i[15]),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(net89),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_3324_),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(net683),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_3360_),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net750),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(net654),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_3343_),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(wbs_dat_i[0]),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(net83),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_3309_),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(net664),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_3335_),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(wbs_dat_i[12]),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(net86),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_3321_),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net752),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(net652),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(_3328_),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(net658),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_3357_),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(net655),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(_3345_),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(net682),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_3340_),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(wbs_dat_i[6]),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(net95),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net738),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_3351_),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(wbs_dat_i[5]),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(net94),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_3333_),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(wbs_dat_i[1]),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(net90),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_3346_),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(net676),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_3329_),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(wbs_dat_i[4]),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net740),
    .X(net312));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold180 (.A(net93),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_3313_),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(net671),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(_3315_),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(net674),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_3314_),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(wbs_dat_i[2]),
    .X(net480));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold187 (.A(net91),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_3330_),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(net680),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net742),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_3350_),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(net653),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_3310_),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(wbs_dat_i[13]),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(net87),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_3341_),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(net689),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_3349_),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(net690),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_3322_),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net716),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net744),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(net675),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_3332_),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(net663),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(_3334_),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(net673),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_3311_),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(wbs_dat_i[3]),
    .X(net500));
 sky130_fd_sc_hd__buf_1 hold207 (.A(net92),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_3331_),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(net677),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net778),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_3347_),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(wbs_dat_i[14]),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(net88),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_3342_),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(net693),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_3348_),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(net695),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_3323_),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(net669),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_3312_),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net780),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(net702),
    .X(net514));
 sky130_fd_sc_hd__buf_1 hold221 (.A(net98),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(_3354_),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(net667),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_3358_),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(net650),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_3359_),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(net649),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(net661),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\mul_wb.p[10] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net758),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_0219_),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\mul_wb.p[9] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_0218_),
    .X(net526));
 sky130_fd_sc_hd__buf_1 hold233 (.A(\mul_wb.p[12] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_0221_),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\mul_wb.p[6] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_0215_),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\mul_wb.p[3] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_0212_),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\mul_wb.p[5] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net760),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_0214_),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\mul_wb.p[4] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(_0213_),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\mul_wb.p[8] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(_0217_),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\mul_wb.p[11] ),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(_0220_),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\mul_wb.p[2] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_0211_),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\mul_wb.p[0] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net746),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_0209_),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\mul_wb.p[1] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_0210_),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\mul_wb.p[7] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_0216_),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(net902),
    .X(net549));
 sky130_fd_sc_hd__buf_12 hold256 (.A(net550),
    .X(la_data_out[0]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(net904),
    .X(net551));
 sky130_fd_sc_hd__buf_12 hold258 (.A(net552),
    .X(la_data_out[7]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(net906),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net748),
    .X(net320));
 sky130_fd_sc_hd__buf_12 hold260 (.A(net554),
    .X(la_data_out[6]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(net908),
    .X(net555));
 sky130_fd_sc_hd__buf_12 hold262 (.A(net556),
    .X(la_data_out[1]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(net910),
    .X(net557));
 sky130_fd_sc_hd__buf_12 hold264 (.A(net558),
    .X(la_data_out[4]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(net912),
    .X(net559));
 sky130_fd_sc_hd__buf_12 hold266 (.A(net560),
    .X(la_data_out[5]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(net914),
    .X(net561));
 sky130_fd_sc_hd__buf_12 hold268 (.A(net562),
    .X(la_data_out[3]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(net916),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net782),
    .X(net321));
 sky130_fd_sc_hd__buf_12 hold270 (.A(net564),
    .X(la_data_out[2]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(net926),
    .X(net565));
 sky130_fd_sc_hd__buf_12 hold272 (.A(net566),
    .X(la_data_out[30]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(net918),
    .X(net567));
 sky130_fd_sc_hd__buf_12 hold274 (.A(net568),
    .X(la_data_out[21]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(net920),
    .X(net569));
 sky130_fd_sc_hd__buf_12 hold276 (.A(net570),
    .X(la_data_out[19]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(net922),
    .X(net571));
 sky130_fd_sc_hd__buf_12 hold278 (.A(net572),
    .X(la_data_out[10]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(net924),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net784),
    .X(net322));
 sky130_fd_sc_hd__buf_12 hold280 (.A(net574),
    .X(la_data_out[9]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(net928),
    .X(net575));
 sky130_fd_sc_hd__buf_12 hold282 (.A(net576),
    .X(la_data_out[13]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(net930),
    .X(net577));
 sky130_fd_sc_hd__buf_12 hold284 (.A(net578),
    .X(la_data_out[18]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(net936),
    .X(net579));
 sky130_fd_sc_hd__buf_12 hold286 (.A(net580),
    .X(la_data_out[26]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(net932),
    .X(net581));
 sky130_fd_sc_hd__buf_12 hold288 (.A(net582),
    .X(la_data_out[8]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(net934),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net718),
    .X(net323));
 sky130_fd_sc_hd__buf_12 hold290 (.A(net584),
    .X(la_data_out[27]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(net944),
    .X(net585));
 sky130_fd_sc_hd__buf_12 hold292 (.A(net586),
    .X(la_data_out[14]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(net938),
    .X(net587));
 sky130_fd_sc_hd__buf_12 hold294 (.A(net588),
    .X(la_data_out[20]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(net942),
    .X(net589));
 sky130_fd_sc_hd__buf_12 hold296 (.A(net590),
    .X(la_data_out[12]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(net940),
    .X(net591));
 sky130_fd_sc_hd__buf_12 hold298 (.A(net592),
    .X(la_data_out[15]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(net946),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net710),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net720),
    .X(net324));
 sky130_fd_sc_hd__buf_12 hold300 (.A(net594),
    .X(la_data_out[16]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(net948),
    .X(net595));
 sky130_fd_sc_hd__buf_12 hold302 (.A(net596),
    .X(la_data_out[22]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(net950),
    .X(net597));
 sky130_fd_sc_hd__buf_12 hold304 (.A(net598),
    .X(la_data_out[29]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(net952),
    .X(net599));
 sky130_fd_sc_hd__buf_12 hold306 (.A(net600),
    .X(la_data_out[23]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(net954),
    .X(net601));
 sky130_fd_sc_hd__buf_12 hold308 (.A(net602),
    .X(la_data_out[31]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(net956),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net730),
    .X(net325));
 sky130_fd_sc_hd__buf_12 hold310 (.A(net604),
    .X(la_data_out[24]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(net958),
    .X(net605));
 sky130_fd_sc_hd__buf_12 hold312 (.A(net606),
    .X(la_data_out[25]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(net960),
    .X(net607));
 sky130_fd_sc_hd__buf_12 hold314 (.A(net608),
    .X(la_data_out[11]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(net962),
    .X(net609));
 sky130_fd_sc_hd__buf_12 hold316 (.A(net610),
    .X(la_data_out[28]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(net964),
    .X(net611));
 sky130_fd_sc_hd__buf_12 hold318 (.A(net612),
    .X(la_data_out[17]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\mul_wb.p[30] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net732),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(_0239_),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\mul_wb.p[29] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(_0238_),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\mul_wb.p[13] ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(_0222_),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\mul_wb.p[14] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(_0223_),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\mul_wb.p[15] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(_0224_),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\mul_wb.p[16] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net726),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(_0225_),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\mul_wb.p[18] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(_0227_),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\mul_wb.p[19] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(_0228_),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\mul_wb.p[17] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(_0226_),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\mul_wb.p[21] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(_0230_),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\mul_wb.p[24] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net728),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(_0233_),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\mul_wb.p[22] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(_0231_),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\mul_wb.p[23] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_0232_),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\mul_wb.p[26] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(_0235_),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\mul_wb.p[20] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(_0229_),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\mul_wb.p[28] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net754),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_0237_),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\mul_wb.p[25] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_0234_),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\mul_wb.p[27] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_0236_),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\mul_wb.b[9] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\mul_wb.a[14] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\mul_wb.a[8] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\mul_wb.b[0] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\mul_wb.l[1] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net756),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\mul_wb.b[15] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\mul_wb.a[0] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(net972),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(net973),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\mul_wb.a[12] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(net976),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(net974),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\mul_wb.l[9] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(net975),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\mul_wb.b[6] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net810),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\mul_wb.b[7] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(net978),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(net977),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\mul_wb.a[13] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(net982),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\mul_wb.l[3] ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(net980),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\mul_wb.l[6] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(net984),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\mul_wb.l[2] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net812),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\mul_wb.l[5] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\mul_wb.b[4] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\mul_wb.b[1] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\mul_wb.a[2] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(net979),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\mul_wb.l[7] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\mul_wb.a[5] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\mul_wb.l[10] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\mul_wb.b[12] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\mul_wb.a[15] ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net802),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\mul_wb.l[8] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(net986),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(net985),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(net983),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(net981),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\mul_wb.a[4] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\mul_wb.l[13] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(net987),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(net989),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\mul_wb.a[3] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net712),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net804),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(net990),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\mul_wb.l[14] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(net988),
    .X(net696));
 sky130_fd_sc_hd__buf_1 hold403 (.A(\mul_wb.reg_b0[15] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(_3619_),
    .X(net698));
 sky130_fd_sc_hd__buf_2 hold405 (.A(\mul_la.reg_b0[15] ),
    .X(net699));
 sky130_fd_sc_hd__buf_2 hold406 (.A(_1808_),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\mul_wb.lob_4.L[15] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(wbs_dat_i[9]),
    .X(net702));
 sky130_fd_sc_hd__clkbuf_2 hold409 (.A(\mul_wb.reg_a0[15] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net766),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_2 hold410 (.A(\mul_la.reg_a0[15] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\mul_wb.lob_4.B[0] ),
    .X(net705));
 sky130_fd_sc_hd__buf_1 hold412 (.A(\mul_wb.reg_a0[14] ),
    .X(net706));
 sky130_fd_sc_hd__buf_1 hold413 (.A(\mul_la.reg_b0[14] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\mul_la.reg_p[30] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\mul_la.lob_4.A[0] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(la_data_in[35]),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(net297),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(net29),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(net298),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net768),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(la_data_in[41]),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(net295),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(net36),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(net296),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(la_data_in[38]),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(net323),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(net32),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(net324),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(la_data_in[10]),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(net299),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net774),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(net2),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(net300),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(la_data_in[37]),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(net327),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(net31),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(net328),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(la_data_in[43]),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(net325),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(net38),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(net326),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net776),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(la_data_in[39]),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(net303),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(net33),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(net304),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(la_data_in[12]),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(net311),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(net4),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(net312),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(la_data_in[36]),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(net313),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net806),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(net30),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(net314),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(la_data_in[46]),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(net319),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(net41),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(net320),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(la_data_in[34]),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(net309),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(net28),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(net310),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net808),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(la_data_in[9]),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(net329),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(net48),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(net330),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(la_data_in[40]),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(net317),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(net35),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(net318),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(la_data_in[8]),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(net301),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net794),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(net47),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(net302),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(la_data_in[18]),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(net335),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(net10),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(net336),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(la_data_in[20]),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(net307),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(net13),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(net308),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net796),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(la_data_in[13]),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(net337),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(net5),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(net338),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(la_data_in[14]),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(net315),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(net6),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(net316),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(la_data_in[15]),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(net321),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net850),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(net7),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(net322),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(la_data_in[42]),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(net355),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(net37),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(net356),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(la_data_in[17]),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(net345),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(net9),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(net346),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net722),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net852),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(la_data_in[27]),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(net341),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(net20),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(net342),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(la_data_in[11]),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(net305),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(net3),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(net306),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(la_data_in[47]),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(net333),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net790),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(net42),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(net334),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(la_data_in[26]),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(net339),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(net19),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(net340),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(la_data_in[32]),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(net331),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(net26),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(net332),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net792),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(la_data_in[19]),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(net369),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(net11),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(net370),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(la_data_in[23]),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(net353),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(net16),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(net354),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(la_data_in[24]),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(net347),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net822),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(net17),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(net348),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(la_data_in[25]),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(net351),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(net18),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(net352),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(la_data_in[31]),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(net349),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(net25),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(net350),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net824),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(la_data_in[29]),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(net357),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(net22),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(net358),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(la_data_in[45]),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(net363),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(net40),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(net364),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(la_data_in[22]),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(net365),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net830),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(net15),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(net366),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(la_data_in[44]),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(net361),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(net39),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(net362),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(la_data_in[30]),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(net343),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(net24),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(net344),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net832),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(la_data_in[28]),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(net367),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(net21),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(net368),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(la_data_in[21]),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(net359),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(net14),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(net360),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(la_data_in[16]),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(net379),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net826),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(net8),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(net380),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(la_data_in[4]),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(net373),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(net43),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(net374),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(la_data_in[6]),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(net375),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(net45),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(net376),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net828),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(la_data_in[33]),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(net371),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(net27),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(net372),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(la_data_in[7]),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(net377),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(net46),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(net378),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(la_data_in[5]),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(net381),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net818),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(net44),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(net382),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(la_data_in[1]),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(net383),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(net12),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(net384),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(la_data_in[3]),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(net385),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(net34),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(net386),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net724),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net820),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(la_data_in[0]),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(net389),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(net1),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(net390),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(la_data_in[2]),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(net387),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(net23),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(net388),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(net101),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(net549),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net786),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(net130),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(net551),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(net129),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(net553),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(net112),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(net555),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(net127),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(net557),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(net128),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(net559),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net788),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(net126),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(net561),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(net123),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(net563),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(net114),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(net567),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(net111),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(net569),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(net102),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(net571),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net834),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(net132),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(net573),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(net124),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(net565),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(net105),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(net575),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(net110),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(net577),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(net131),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(net581),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net836),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(net120),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(net583),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(net119),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(net579),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(net113),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(net587),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(net107),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(net591),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(net104),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(net589),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net858),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(net106),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(net585),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(net108),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(net593),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(net115),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(net595),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(net122),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(net597),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(net116),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(net599),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net860),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(net125),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(net601),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(net117),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(net603),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(net118),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(net605),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(net103),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(net607),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(net121),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(net609),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net846),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(net109),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(net611),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(wbs_adr_i[22]),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(_3297_),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(_3303_),
    .X(net968));
 sky130_fd_sc_hd__buf_1 hold675 (.A(\mul_wb.reg_b0[14] ),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(_3498_),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(\mul_wb.b[10] ),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\mul_wb.l[4] ),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net848),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\mul_wb.b[5] ),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\mul_wb.l[12] ),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\mul_wb.b[8] ),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\mul_wb.a[1] ),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(\mul_wb.a[9] ),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\mul_wb.a[7] ),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(\mul_wb.a[6] ),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\mul_wb.b[13] ),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(\mul_wb.b[3] ),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\mul_wb.b[2] ),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net838),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\mul_wb.l[0] ),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\mul_wb.b[14] ),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(\mul_wb.b[11] ),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\mul_wb.l[11] ),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\mul_wb.a[11] ),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\mul_wb.l[15] ),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\mul_wb.a[10] ),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(\mul_wb.p[31] ),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\mul_wb.reg_a0[12] ),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(_3392_),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net762),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net840),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(_3393_),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net842),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net844),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net854),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net856),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net814),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net816),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net874),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net876),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net866),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net764),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net868),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net870),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net872),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net878),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net880),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net862),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net864),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net882),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net884),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net886),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net734),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(net888),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net890),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net892),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net898),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net900),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(net894),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net896),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(wbs_adr_i[1]),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net61),
    .X(net392));
 sky130_fd_sc_hd__buf_1 hold99 (.A(_3304_),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(net895),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(net767),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input100 (.A(wbs_we_i),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(net815),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(net887),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(net771),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(net859),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(net843),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(net819),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(net823),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(net827),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(net807),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(net723),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(net795),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(net855),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(net835),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(net899),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(net851),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(net831),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(net811),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(net875),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(net751),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(net711),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(net799),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(net743),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(net727),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(net719),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(net735),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(net891),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(net759),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(net715),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(net787),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(net731),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(net847),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input4 (.A(net739),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(net839),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(net747),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(net803),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(net867),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(net883),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(net871),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(net879),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(net763),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(net755),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(wb_rst_i),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input5 (.A(net775),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(net410),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(wbs_adr_i[10]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(wbs_adr_i[11]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(wbs_adr_i[12]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(wbs_adr_i[13]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(wbs_adr_i[14]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(wbs_adr_i[15]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(wbs_adr_i[16]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(wbs_adr_i[17]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(wbs_adr_i[18]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(net779),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(wbs_adr_i[19]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(net391),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(wbs_adr_i[20]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(wbs_adr_i[21]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(net966),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(wbs_adr_i[23]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(wbs_adr_i[24]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(wbs_adr_i[25]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(net426),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(wbs_adr_i[27]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input7 (.A(net783),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(wbs_adr_i[28]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(wbs_adr_i[29]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(net404),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(wbs_adr_i[30]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(wbs_adr_i[31]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(net395),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(wbs_adr_i[4]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(wbs_adr_i[5]),
    .X(net77));
 sky130_fd_sc_hd__buf_1 input78 (.A(wbs_adr_i[6]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(wbs_adr_i[7]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(net863),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input80 (.A(wbs_adr_i[8]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(wbs_adr_i[9]),
    .X(net81));
 sky130_fd_sc_hd__dlymetal6s2s_1 input82 (.A(wbs_cyc_i),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(net446),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(net420),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(net400),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(net451),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(net487),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(net505),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(net439),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(net791),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(net468),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(net480),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(net500),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input93 (.A(net473),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(net465),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(net462),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(net432),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(net414),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(net514),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(wbs_stb_i),
    .X(net99));
 sky130_fd_sc_hd__buf_1 max_cap166 (.A(_2042_),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_4 max_cap180 (.A(_2142_),
    .X(net180));
 sky130_fd_sc_hd__buf_2 max_cap184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 max_cap185 (.A(_1967_),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_4 max_cap205 (.A(_3773_),
    .X(net205));
 sky130_fd_sc_hd__buf_4 max_cap211 (.A(_3613_),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 max_cap215 (.A(_2060_),
    .X(net215));
 sky130_fd_sc_hd__buf_6 max_cap226 (.A(_1696_),
    .X(net226));
 sky130_fd_sc_hd__buf_1 max_cap231 (.A(_1799_),
    .X(net231));
 sky130_fd_sc_hd__buf_2 max_cap234 (.A(_1646_),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_2 max_cap238 (.A(_3545_),
    .X(net238));
 sky130_fd_sc_hd__buf_1 max_cap240 (.A(_3530_),
    .X(net240));
 sky130_fd_sc_hd__buf_2 max_cap241 (.A(_3444_),
    .X(net241));
 sky130_fd_sc_hd__buf_4 max_cap242 (.A(_3498_),
    .X(net242));
 sky130_fd_sc_hd__buf_6 max_cap245 (.A(_3483_),
    .X(net245));
 sky130_fd_sc_hd__buf_4 max_cap247 (.A(_3397_),
    .X(net247));
 sky130_fd_sc_hd__buf_6 output101 (.A(net903),
    .X(net550));
 sky130_fd_sc_hd__buf_6 output102 (.A(net923),
    .X(net572));
 sky130_fd_sc_hd__buf_6 output103 (.A(net961),
    .X(net608));
 sky130_fd_sc_hd__buf_6 output104 (.A(net943),
    .X(net590));
 sky130_fd_sc_hd__buf_6 output105 (.A(net929),
    .X(net576));
 sky130_fd_sc_hd__buf_6 output106 (.A(net945),
    .X(net586));
 sky130_fd_sc_hd__buf_6 output107 (.A(net941),
    .X(net592));
 sky130_fd_sc_hd__buf_6 output108 (.A(net947),
    .X(net594));
 sky130_fd_sc_hd__buf_6 output109 (.A(net965),
    .X(net612));
 sky130_fd_sc_hd__buf_6 output110 (.A(net931),
    .X(net578));
 sky130_fd_sc_hd__buf_6 output111 (.A(net921),
    .X(net570));
 sky130_fd_sc_hd__buf_6 output112 (.A(net909),
    .X(net556));
 sky130_fd_sc_hd__buf_6 output113 (.A(net939),
    .X(net588));
 sky130_fd_sc_hd__buf_6 output114 (.A(net919),
    .X(net568));
 sky130_fd_sc_hd__buf_6 output115 (.A(net949),
    .X(net596));
 sky130_fd_sc_hd__buf_6 output116 (.A(net953),
    .X(net600));
 sky130_fd_sc_hd__buf_6 output117 (.A(net957),
    .X(net604));
 sky130_fd_sc_hd__buf_6 output118 (.A(net959),
    .X(net606));
 sky130_fd_sc_hd__buf_6 output119 (.A(net937),
    .X(net580));
 sky130_fd_sc_hd__buf_6 output120 (.A(net935),
    .X(net584));
 sky130_fd_sc_hd__buf_6 output121 (.A(net963),
    .X(net610));
 sky130_fd_sc_hd__buf_6 output122 (.A(net951),
    .X(net598));
 sky130_fd_sc_hd__buf_6 output123 (.A(net917),
    .X(net564));
 sky130_fd_sc_hd__buf_6 output124 (.A(net927),
    .X(net566));
 sky130_fd_sc_hd__buf_6 output125 (.A(net955),
    .X(net602));
 sky130_fd_sc_hd__buf_6 output126 (.A(net915),
    .X(net562));
 sky130_fd_sc_hd__buf_6 output127 (.A(net911),
    .X(net558));
 sky130_fd_sc_hd__buf_6 output128 (.A(net913),
    .X(net560));
 sky130_fd_sc_hd__buf_6 output129 (.A(net907),
    .X(net554));
 sky130_fd_sc_hd__buf_6 output130 (.A(net905),
    .X(net552));
 sky130_fd_sc_hd__buf_6 output131 (.A(net933),
    .X(net582));
 sky130_fd_sc_hd__buf_6 output132 (.A(net925),
    .X(net574));
 sky130_fd_sc_hd__buf_12 output133 (.A(net133),
    .X(wbs_ack_o));
 sky130_fd_sc_hd__buf_12 output134 (.A(net134),
    .X(wbs_dat_o[0]));
 sky130_fd_sc_hd__buf_12 output135 (.A(net135),
    .X(wbs_dat_o[10]));
 sky130_fd_sc_hd__buf_12 output136 (.A(net136),
    .X(wbs_dat_o[11]));
 sky130_fd_sc_hd__buf_12 output137 (.A(net137),
    .X(wbs_dat_o[12]));
 sky130_fd_sc_hd__buf_12 output138 (.A(net138),
    .X(wbs_dat_o[13]));
 sky130_fd_sc_hd__buf_12 output139 (.A(net139),
    .X(wbs_dat_o[14]));
 sky130_fd_sc_hd__buf_12 output140 (.A(net140),
    .X(wbs_dat_o[15]));
 sky130_fd_sc_hd__buf_12 output141 (.A(net141),
    .X(wbs_dat_o[16]));
 sky130_fd_sc_hd__buf_12 output142 (.A(net142),
    .X(wbs_dat_o[17]));
 sky130_fd_sc_hd__buf_12 output143 (.A(net143),
    .X(wbs_dat_o[18]));
 sky130_fd_sc_hd__buf_12 output144 (.A(net144),
    .X(wbs_dat_o[19]));
 sky130_fd_sc_hd__buf_12 output145 (.A(net145),
    .X(wbs_dat_o[1]));
 sky130_fd_sc_hd__buf_12 output146 (.A(net146),
    .X(wbs_dat_o[20]));
 sky130_fd_sc_hd__buf_12 output147 (.A(net147),
    .X(wbs_dat_o[21]));
 sky130_fd_sc_hd__buf_12 output148 (.A(net148),
    .X(wbs_dat_o[22]));
 sky130_fd_sc_hd__buf_12 output149 (.A(net149),
    .X(wbs_dat_o[23]));
 sky130_fd_sc_hd__buf_12 output150 (.A(net150),
    .X(wbs_dat_o[24]));
 sky130_fd_sc_hd__buf_12 output151 (.A(net151),
    .X(wbs_dat_o[25]));
 sky130_fd_sc_hd__buf_12 output152 (.A(net152),
    .X(wbs_dat_o[26]));
 sky130_fd_sc_hd__buf_12 output153 (.A(net153),
    .X(wbs_dat_o[27]));
 sky130_fd_sc_hd__buf_12 output154 (.A(net154),
    .X(wbs_dat_o[28]));
 sky130_fd_sc_hd__buf_12 output155 (.A(net155),
    .X(wbs_dat_o[29]));
 sky130_fd_sc_hd__buf_12 output156 (.A(net156),
    .X(wbs_dat_o[2]));
 sky130_fd_sc_hd__buf_12 output157 (.A(net157),
    .X(wbs_dat_o[30]));
 sky130_fd_sc_hd__buf_12 output158 (.A(net158),
    .X(wbs_dat_o[31]));
 sky130_fd_sc_hd__buf_12 output159 (.A(net159),
    .X(wbs_dat_o[3]));
 sky130_fd_sc_hd__buf_12 output160 (.A(net160),
    .X(wbs_dat_o[4]));
 sky130_fd_sc_hd__buf_12 output161 (.A(net161),
    .X(wbs_dat_o[5]));
 sky130_fd_sc_hd__buf_12 output162 (.A(net162),
    .X(wbs_dat_o[6]));
 sky130_fd_sc_hd__buf_12 output163 (.A(net163),
    .X(wbs_dat_o[7]));
 sky130_fd_sc_hd__buf_12 output164 (.A(net164),
    .X(wbs_dat_o[8]));
 sky130_fd_sc_hd__buf_12 output165 (.A(net165),
    .X(wbs_dat_o[9]));
 sky130_fd_sc_hd__conb_1 wb_RAxM_294 (.LO(net294));
 sky130_fd_sc_hd__clkbuf_4 wire171 (.A(_1847_),
    .X(net171));
 sky130_fd_sc_hd__buf_4 wire212 (.A(_3608_),
    .X(net212));
 sky130_fd_sc_hd__buf_1 wire228 (.A(_3473_),
    .X(net228));
 sky130_fd_sc_hd__buf_2 wire239 (.A(_3543_),
    .X(net239));
 assign wbs_sta_o = net294;
endmodule

