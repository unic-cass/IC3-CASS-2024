VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 17.720 500.000 18.320 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 87.080 500.000 87.680 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 156.440 500.000 157.040 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 225.800 500.000 226.400 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 295.160 500.000 295.760 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 364.520 500.000 365.120 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 433.880 500.000 434.480 ;
    END
  END io_in[6]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 63.960 500.000 64.560 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 133.320 500.000 133.920 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 202.680 500.000 203.280 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 272.040 500.000 272.640 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 341.400 500.000 342.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 410.760 500.000 411.360 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 480.120 500.000 480.720 ;
    END
  END io_oeb[6]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 40.840 500.000 41.440 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 110.200 500.000 110.800 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 179.560 500.000 180.160 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 248.920 500.000 249.520 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 318.280 500.000 318.880 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 387.640 500.000 388.240 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 457.000 500.000 457.600 ;
    END
  END io_out[6]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END wb_clk_i
  OBS
      LAYER nwell ;
        RECT 5.330 485.465 494.230 487.070 ;
        RECT 5.330 480.025 494.230 482.855 ;
        RECT 5.330 474.585 494.230 477.415 ;
        RECT 5.330 469.145 494.230 471.975 ;
        RECT 5.330 463.705 494.230 466.535 ;
        RECT 5.330 458.265 494.230 461.095 ;
        RECT 5.330 452.825 494.230 455.655 ;
        RECT 5.330 447.385 494.230 450.215 ;
        RECT 5.330 441.945 494.230 444.775 ;
        RECT 5.330 436.505 494.230 439.335 ;
        RECT 5.330 431.065 494.230 433.895 ;
        RECT 5.330 425.625 494.230 428.455 ;
        RECT 5.330 420.185 494.230 423.015 ;
        RECT 5.330 414.745 494.230 417.575 ;
        RECT 5.330 409.305 494.230 412.135 ;
        RECT 5.330 403.865 494.230 406.695 ;
        RECT 5.330 398.425 494.230 401.255 ;
        RECT 5.330 392.985 494.230 395.815 ;
        RECT 5.330 387.545 494.230 390.375 ;
        RECT 5.330 382.105 494.230 384.935 ;
        RECT 5.330 376.665 494.230 379.495 ;
        RECT 5.330 371.225 494.230 374.055 ;
        RECT 5.330 365.785 494.230 368.615 ;
        RECT 5.330 360.345 494.230 363.175 ;
        RECT 5.330 354.905 494.230 357.735 ;
        RECT 5.330 349.465 494.230 352.295 ;
        RECT 5.330 344.025 494.230 346.855 ;
        RECT 5.330 338.585 494.230 341.415 ;
        RECT 5.330 333.145 494.230 335.975 ;
        RECT 5.330 327.705 494.230 330.535 ;
        RECT 5.330 322.265 494.230 325.095 ;
        RECT 5.330 316.825 494.230 319.655 ;
        RECT 5.330 311.385 494.230 314.215 ;
        RECT 5.330 305.945 494.230 308.775 ;
        RECT 5.330 300.505 494.230 303.335 ;
        RECT 5.330 295.065 494.230 297.895 ;
        RECT 5.330 289.625 494.230 292.455 ;
        RECT 5.330 284.185 494.230 287.015 ;
        RECT 5.330 278.745 494.230 281.575 ;
        RECT 5.330 273.305 494.230 276.135 ;
        RECT 5.330 267.865 494.230 270.695 ;
        RECT 5.330 262.425 494.230 265.255 ;
        RECT 5.330 256.985 494.230 259.815 ;
        RECT 5.330 251.545 494.230 254.375 ;
        RECT 5.330 246.105 494.230 248.935 ;
        RECT 5.330 240.665 494.230 243.495 ;
        RECT 5.330 235.225 494.230 238.055 ;
        RECT 5.330 229.785 494.230 232.615 ;
        RECT 5.330 224.345 494.230 227.175 ;
        RECT 5.330 218.905 494.230 221.735 ;
        RECT 5.330 213.465 494.230 216.295 ;
        RECT 5.330 208.025 494.230 210.855 ;
        RECT 5.330 202.585 494.230 205.415 ;
        RECT 5.330 197.145 494.230 199.975 ;
        RECT 5.330 191.705 494.230 194.535 ;
        RECT 5.330 186.265 494.230 189.095 ;
        RECT 5.330 180.825 494.230 183.655 ;
        RECT 5.330 175.385 494.230 178.215 ;
        RECT 5.330 169.945 494.230 172.775 ;
        RECT 5.330 164.505 494.230 167.335 ;
        RECT 5.330 159.065 494.230 161.895 ;
        RECT 5.330 153.625 494.230 156.455 ;
        RECT 5.330 148.185 494.230 151.015 ;
        RECT 5.330 142.745 494.230 145.575 ;
        RECT 5.330 137.305 494.230 140.135 ;
        RECT 5.330 131.865 494.230 134.695 ;
        RECT 5.330 126.425 494.230 129.255 ;
        RECT 5.330 120.985 494.230 123.815 ;
        RECT 5.330 115.545 494.230 118.375 ;
        RECT 5.330 110.105 494.230 112.935 ;
        RECT 5.330 104.665 494.230 107.495 ;
        RECT 5.330 99.225 494.230 102.055 ;
        RECT 5.330 93.785 494.230 96.615 ;
        RECT 5.330 88.345 494.230 91.175 ;
        RECT 5.330 82.905 494.230 85.735 ;
        RECT 5.330 77.465 494.230 80.295 ;
        RECT 5.330 72.025 494.230 74.855 ;
        RECT 5.330 66.585 494.230 69.415 ;
        RECT 5.330 61.145 494.230 63.975 ;
        RECT 5.330 55.705 494.230 58.535 ;
        RECT 5.330 50.265 494.230 53.095 ;
        RECT 5.330 44.825 494.230 47.655 ;
        RECT 5.330 39.385 494.230 42.215 ;
        RECT 5.330 33.945 494.230 36.775 ;
        RECT 5.330 28.505 494.230 31.335 ;
        RECT 5.330 23.065 494.230 25.895 ;
        RECT 5.330 17.625 494.230 20.455 ;
        RECT 5.330 12.185 494.230 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 5.520 10.640 494.430 487.120 ;
      LAYER met2 ;
        RECT 21.070 4.280 494.410 487.065 ;
        RECT 21.070 4.000 249.590 4.280 ;
        RECT 250.430 4.000 494.410 4.280 ;
      LAYER met3 ;
        RECT 21.050 481.120 496.000 487.045 ;
        RECT 21.050 479.720 495.600 481.120 ;
        RECT 21.050 458.000 496.000 479.720 ;
        RECT 21.050 456.600 495.600 458.000 ;
        RECT 21.050 434.880 496.000 456.600 ;
        RECT 21.050 433.480 495.600 434.880 ;
        RECT 21.050 411.760 496.000 433.480 ;
        RECT 21.050 410.360 495.600 411.760 ;
        RECT 21.050 388.640 496.000 410.360 ;
        RECT 21.050 387.240 495.600 388.640 ;
        RECT 21.050 365.520 496.000 387.240 ;
        RECT 21.050 364.120 495.600 365.520 ;
        RECT 21.050 342.400 496.000 364.120 ;
        RECT 21.050 341.000 495.600 342.400 ;
        RECT 21.050 319.280 496.000 341.000 ;
        RECT 21.050 317.880 495.600 319.280 ;
        RECT 21.050 296.160 496.000 317.880 ;
        RECT 21.050 294.760 495.600 296.160 ;
        RECT 21.050 273.040 496.000 294.760 ;
        RECT 21.050 271.640 495.600 273.040 ;
        RECT 21.050 249.920 496.000 271.640 ;
        RECT 21.050 248.520 495.600 249.920 ;
        RECT 21.050 226.800 496.000 248.520 ;
        RECT 21.050 225.400 495.600 226.800 ;
        RECT 21.050 203.680 496.000 225.400 ;
        RECT 21.050 202.280 495.600 203.680 ;
        RECT 21.050 180.560 496.000 202.280 ;
        RECT 21.050 179.160 495.600 180.560 ;
        RECT 21.050 157.440 496.000 179.160 ;
        RECT 21.050 156.040 495.600 157.440 ;
        RECT 21.050 134.320 496.000 156.040 ;
        RECT 21.050 132.920 495.600 134.320 ;
        RECT 21.050 111.200 496.000 132.920 ;
        RECT 21.050 109.800 495.600 111.200 ;
        RECT 21.050 88.080 496.000 109.800 ;
        RECT 21.050 86.680 495.600 88.080 ;
        RECT 21.050 64.960 496.000 86.680 ;
        RECT 21.050 63.560 495.600 64.960 ;
        RECT 21.050 41.840 496.000 63.560 ;
        RECT 21.050 40.440 495.600 41.840 ;
        RECT 21.050 18.720 496.000 40.440 ;
        RECT 21.050 17.320 495.600 18.720 ;
        RECT 21.050 10.715 496.000 17.320 ;
  END
END user_proj_example
END LIBRARY

