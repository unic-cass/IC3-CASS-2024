VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_RAxM
  CLASS BLOCK ;
  FOREIGN wb_RAxM ;
  ORIGIN 0.000 0.000 ;
  SIZE 324.040 BY 334.760 ;
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 5.480 324.040 6.080 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 320.040 46.280 324.040 46.880 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 50.360 324.040 50.960 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 54.440 324.040 55.040 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 58.520 324.040 59.120 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 62.600 324.040 63.200 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 66.680 324.040 67.280 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 70.760 324.040 71.360 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 74.840 324.040 75.440 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 78.920 324.040 79.520 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 83.000 324.040 83.600 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 9.560 324.040 10.160 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 87.080 324.040 87.680 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 91.160 324.040 91.760 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 95.240 324.040 95.840 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 99.320 324.040 99.920 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 103.400 324.040 104.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 107.480 324.040 108.080 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 111.560 324.040 112.160 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 115.640 324.040 116.240 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 119.720 324.040 120.320 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 123.800 324.040 124.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 13.640 324.040 14.240 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 127.880 324.040 128.480 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 131.960 324.040 132.560 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 136.040 324.040 136.640 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 140.120 324.040 140.720 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 144.200 324.040 144.800 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 148.280 324.040 148.880 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 152.360 324.040 152.960 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 156.440 324.040 157.040 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 160.520 324.040 161.120 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 164.600 324.040 165.200 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 320.040 17.720 324.040 18.320 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 168.680 324.040 169.280 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 172.760 324.040 173.360 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 176.840 324.040 177.440 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 180.920 324.040 181.520 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 185.000 324.040 185.600 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 189.080 324.040 189.680 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 193.160 324.040 193.760 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 197.240 324.040 197.840 ;
    END
  END la_data_in[47]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 21.800 324.040 22.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 25.880 324.040 26.480 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 320.040 29.960 324.040 30.560 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 34.040 324.040 34.640 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 38.120 324.040 38.720 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 320.040 42.200 324.040 42.800 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 201.320 324.040 201.920 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 242.120 324.040 242.720 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 246.200 324.040 246.800 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 250.280 324.040 250.880 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 254.360 324.040 254.960 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 258.440 324.040 259.040 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 262.520 324.040 263.120 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 266.600 324.040 267.200 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 270.680 324.040 271.280 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 274.760 324.040 275.360 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 278.840 324.040 279.440 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 205.400 324.040 206.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 282.920 324.040 283.520 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 287.000 324.040 287.600 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 291.080 324.040 291.680 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 295.160 324.040 295.760 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 299.240 324.040 299.840 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 303.320 324.040 303.920 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 307.400 324.040 308.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 311.480 324.040 312.080 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 315.560 324.040 316.160 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 319.640 324.040 320.240 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 209.480 324.040 210.080 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 323.720 324.040 324.320 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 327.800 324.040 328.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 213.560 324.040 214.160 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 217.640 324.040 218.240 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 221.720 324.040 222.320 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 225.800 324.040 226.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 229.880 324.040 230.480 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 233.960 324.040 234.560 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 320.040 238.040 324.040 238.640 ;
    END
  END la_data_out[9]
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 323.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 323.920 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 323.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 323.920 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 252.630 0.000 252.910 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 277.470 0.000 277.750 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sta_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END wbs_sta_o
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER nwell ;
        RECT 5.330 322.265 318.510 323.870 ;
        RECT 5.330 316.825 318.510 319.655 ;
        RECT 5.330 311.385 318.510 314.215 ;
        RECT 5.330 305.945 318.510 308.775 ;
        RECT 5.330 300.505 318.510 303.335 ;
        RECT 5.330 295.065 318.510 297.895 ;
        RECT 5.330 289.625 318.510 292.455 ;
        RECT 5.330 284.185 318.510 287.015 ;
        RECT 5.330 278.745 318.510 281.575 ;
        RECT 5.330 273.305 318.510 276.135 ;
        RECT 5.330 267.865 318.510 270.695 ;
        RECT 5.330 262.425 318.510 265.255 ;
        RECT 5.330 256.985 318.510 259.815 ;
        RECT 5.330 251.545 318.510 254.375 ;
        RECT 5.330 246.105 318.510 248.935 ;
        RECT 5.330 240.665 318.510 243.495 ;
        RECT 5.330 235.225 318.510 238.055 ;
        RECT 5.330 229.785 318.510 232.615 ;
        RECT 5.330 224.345 318.510 227.175 ;
        RECT 5.330 218.905 318.510 221.735 ;
        RECT 5.330 213.465 318.510 216.295 ;
        RECT 5.330 208.025 318.510 210.855 ;
        RECT 5.330 202.585 318.510 205.415 ;
        RECT 5.330 197.145 318.510 199.975 ;
        RECT 5.330 191.705 318.510 194.535 ;
        RECT 5.330 186.265 318.510 189.095 ;
        RECT 5.330 180.825 318.510 183.655 ;
        RECT 5.330 175.385 318.510 178.215 ;
        RECT 5.330 169.945 318.510 172.775 ;
        RECT 5.330 164.505 318.510 167.335 ;
        RECT 5.330 159.065 318.510 161.895 ;
        RECT 5.330 153.625 318.510 156.455 ;
        RECT 5.330 148.185 318.510 151.015 ;
        RECT 5.330 142.745 318.510 145.575 ;
        RECT 5.330 137.305 318.510 140.135 ;
        RECT 5.330 131.865 318.510 134.695 ;
        RECT 5.330 126.425 318.510 129.255 ;
        RECT 5.330 120.985 318.510 123.815 ;
        RECT 5.330 115.545 318.510 118.375 ;
        RECT 5.330 110.105 318.510 112.935 ;
        RECT 5.330 104.665 318.510 107.495 ;
        RECT 5.330 99.225 318.510 102.055 ;
        RECT 5.330 93.785 318.510 96.615 ;
        RECT 5.330 88.345 318.510 91.175 ;
        RECT 5.330 82.905 318.510 85.735 ;
        RECT 5.330 77.465 318.510 80.295 ;
        RECT 5.330 72.025 318.510 74.855 ;
        RECT 5.330 66.585 318.510 69.415 ;
        RECT 5.330 61.145 318.510 63.975 ;
        RECT 5.330 55.705 318.510 58.535 ;
        RECT 5.330 50.265 318.510 53.095 ;
        RECT 5.330 44.825 318.510 47.655 ;
        RECT 5.330 39.385 318.510 42.215 ;
        RECT 5.330 33.945 318.510 36.775 ;
        RECT 5.330 28.505 318.510 31.335 ;
        RECT 5.330 23.065 318.510 25.895 ;
        RECT 5.330 17.625 318.510 20.455 ;
        RECT 5.330 12.185 318.510 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 318.320 323.765 ;
      LAYER met1 ;
        RECT 5.520 6.500 321.470 324.660 ;
      LAYER met2 ;
        RECT 5.610 4.280 321.450 328.285 ;
        RECT 5.610 3.670 20.510 4.280 ;
        RECT 21.350 3.670 23.270 4.280 ;
        RECT 24.110 3.670 26.030 4.280 ;
        RECT 26.870 3.670 28.790 4.280 ;
        RECT 29.630 3.670 31.550 4.280 ;
        RECT 32.390 3.670 34.310 4.280 ;
        RECT 35.150 3.670 37.070 4.280 ;
        RECT 37.910 3.670 39.830 4.280 ;
        RECT 40.670 3.670 42.590 4.280 ;
        RECT 43.430 3.670 45.350 4.280 ;
        RECT 46.190 3.670 48.110 4.280 ;
        RECT 48.950 3.670 50.870 4.280 ;
        RECT 51.710 3.670 53.630 4.280 ;
        RECT 54.470 3.670 56.390 4.280 ;
        RECT 57.230 3.670 59.150 4.280 ;
        RECT 59.990 3.670 61.910 4.280 ;
        RECT 62.750 3.670 64.670 4.280 ;
        RECT 65.510 3.670 67.430 4.280 ;
        RECT 68.270 3.670 70.190 4.280 ;
        RECT 71.030 3.670 72.950 4.280 ;
        RECT 73.790 3.670 75.710 4.280 ;
        RECT 76.550 3.670 78.470 4.280 ;
        RECT 79.310 3.670 81.230 4.280 ;
        RECT 82.070 3.670 83.990 4.280 ;
        RECT 84.830 3.670 86.750 4.280 ;
        RECT 87.590 3.670 89.510 4.280 ;
        RECT 90.350 3.670 92.270 4.280 ;
        RECT 93.110 3.670 95.030 4.280 ;
        RECT 95.870 3.670 97.790 4.280 ;
        RECT 98.630 3.670 100.550 4.280 ;
        RECT 101.390 3.670 103.310 4.280 ;
        RECT 104.150 3.670 106.070 4.280 ;
        RECT 106.910 3.670 108.830 4.280 ;
        RECT 109.670 3.670 111.590 4.280 ;
        RECT 112.430 3.670 114.350 4.280 ;
        RECT 115.190 3.670 117.110 4.280 ;
        RECT 117.950 3.670 119.870 4.280 ;
        RECT 120.710 3.670 122.630 4.280 ;
        RECT 123.470 3.670 125.390 4.280 ;
        RECT 126.230 3.670 128.150 4.280 ;
        RECT 128.990 3.670 130.910 4.280 ;
        RECT 131.750 3.670 133.670 4.280 ;
        RECT 134.510 3.670 136.430 4.280 ;
        RECT 137.270 3.670 139.190 4.280 ;
        RECT 140.030 3.670 141.950 4.280 ;
        RECT 142.790 3.670 144.710 4.280 ;
        RECT 145.550 3.670 147.470 4.280 ;
        RECT 148.310 3.670 150.230 4.280 ;
        RECT 151.070 3.670 152.990 4.280 ;
        RECT 153.830 3.670 155.750 4.280 ;
        RECT 156.590 3.670 158.510 4.280 ;
        RECT 159.350 3.670 161.270 4.280 ;
        RECT 162.110 3.670 164.030 4.280 ;
        RECT 164.870 3.670 166.790 4.280 ;
        RECT 167.630 3.670 169.550 4.280 ;
        RECT 170.390 3.670 172.310 4.280 ;
        RECT 173.150 3.670 175.070 4.280 ;
        RECT 175.910 3.670 177.830 4.280 ;
        RECT 178.670 3.670 180.590 4.280 ;
        RECT 181.430 3.670 183.350 4.280 ;
        RECT 184.190 3.670 186.110 4.280 ;
        RECT 186.950 3.670 188.870 4.280 ;
        RECT 189.710 3.670 191.630 4.280 ;
        RECT 192.470 3.670 194.390 4.280 ;
        RECT 195.230 3.670 197.150 4.280 ;
        RECT 197.990 3.670 199.910 4.280 ;
        RECT 200.750 3.670 202.670 4.280 ;
        RECT 203.510 3.670 205.430 4.280 ;
        RECT 206.270 3.670 208.190 4.280 ;
        RECT 209.030 3.670 210.950 4.280 ;
        RECT 211.790 3.670 213.710 4.280 ;
        RECT 214.550 3.670 216.470 4.280 ;
        RECT 217.310 3.670 219.230 4.280 ;
        RECT 220.070 3.670 221.990 4.280 ;
        RECT 222.830 3.670 224.750 4.280 ;
        RECT 225.590 3.670 227.510 4.280 ;
        RECT 228.350 3.670 230.270 4.280 ;
        RECT 231.110 3.670 233.030 4.280 ;
        RECT 233.870 3.670 235.790 4.280 ;
        RECT 236.630 3.670 238.550 4.280 ;
        RECT 239.390 3.670 241.310 4.280 ;
        RECT 242.150 3.670 244.070 4.280 ;
        RECT 244.910 3.670 246.830 4.280 ;
        RECT 247.670 3.670 249.590 4.280 ;
        RECT 250.430 3.670 252.350 4.280 ;
        RECT 253.190 3.670 255.110 4.280 ;
        RECT 255.950 3.670 257.870 4.280 ;
        RECT 258.710 3.670 260.630 4.280 ;
        RECT 261.470 3.670 263.390 4.280 ;
        RECT 264.230 3.670 266.150 4.280 ;
        RECT 266.990 3.670 268.910 4.280 ;
        RECT 269.750 3.670 271.670 4.280 ;
        RECT 272.510 3.670 274.430 4.280 ;
        RECT 275.270 3.670 277.190 4.280 ;
        RECT 278.030 3.670 279.950 4.280 ;
        RECT 280.790 3.670 282.710 4.280 ;
        RECT 283.550 3.670 285.470 4.280 ;
        RECT 286.310 3.670 288.230 4.280 ;
        RECT 289.070 3.670 290.990 4.280 ;
        RECT 291.830 3.670 293.750 4.280 ;
        RECT 294.590 3.670 296.510 4.280 ;
        RECT 297.350 3.670 299.270 4.280 ;
        RECT 300.110 3.670 302.030 4.280 ;
        RECT 302.870 3.670 321.450 4.280 ;
      LAYER met3 ;
        RECT 5.585 327.400 319.640 328.265 ;
        RECT 5.585 324.720 321.475 327.400 ;
        RECT 5.585 323.320 319.640 324.720 ;
        RECT 5.585 320.640 321.475 323.320 ;
        RECT 5.585 319.240 319.640 320.640 ;
        RECT 5.585 316.560 321.475 319.240 ;
        RECT 5.585 315.160 319.640 316.560 ;
        RECT 5.585 312.480 321.475 315.160 ;
        RECT 5.585 311.080 319.640 312.480 ;
        RECT 5.585 308.400 321.475 311.080 ;
        RECT 5.585 307.000 319.640 308.400 ;
        RECT 5.585 304.320 321.475 307.000 ;
        RECT 5.585 302.920 319.640 304.320 ;
        RECT 5.585 300.240 321.475 302.920 ;
        RECT 5.585 298.840 319.640 300.240 ;
        RECT 5.585 296.160 321.475 298.840 ;
        RECT 5.585 294.760 319.640 296.160 ;
        RECT 5.585 292.080 321.475 294.760 ;
        RECT 5.585 290.680 319.640 292.080 ;
        RECT 5.585 288.000 321.475 290.680 ;
        RECT 5.585 286.600 319.640 288.000 ;
        RECT 5.585 283.920 321.475 286.600 ;
        RECT 5.585 282.520 319.640 283.920 ;
        RECT 5.585 279.840 321.475 282.520 ;
        RECT 5.585 278.440 319.640 279.840 ;
        RECT 5.585 275.760 321.475 278.440 ;
        RECT 5.585 274.360 319.640 275.760 ;
        RECT 5.585 271.680 321.475 274.360 ;
        RECT 5.585 270.280 319.640 271.680 ;
        RECT 5.585 267.600 321.475 270.280 ;
        RECT 5.585 266.200 319.640 267.600 ;
        RECT 5.585 263.520 321.475 266.200 ;
        RECT 5.585 262.120 319.640 263.520 ;
        RECT 5.585 259.440 321.475 262.120 ;
        RECT 5.585 258.040 319.640 259.440 ;
        RECT 5.585 255.360 321.475 258.040 ;
        RECT 5.585 253.960 319.640 255.360 ;
        RECT 5.585 251.280 321.475 253.960 ;
        RECT 5.585 249.880 319.640 251.280 ;
        RECT 5.585 247.200 321.475 249.880 ;
        RECT 5.585 245.800 319.640 247.200 ;
        RECT 5.585 243.120 321.475 245.800 ;
        RECT 5.585 241.720 319.640 243.120 ;
        RECT 5.585 239.040 321.475 241.720 ;
        RECT 5.585 237.640 319.640 239.040 ;
        RECT 5.585 234.960 321.475 237.640 ;
        RECT 5.585 233.560 319.640 234.960 ;
        RECT 5.585 230.880 321.475 233.560 ;
        RECT 5.585 229.480 319.640 230.880 ;
        RECT 5.585 226.800 321.475 229.480 ;
        RECT 5.585 225.400 319.640 226.800 ;
        RECT 5.585 222.720 321.475 225.400 ;
        RECT 5.585 221.320 319.640 222.720 ;
        RECT 5.585 218.640 321.475 221.320 ;
        RECT 5.585 217.240 319.640 218.640 ;
        RECT 5.585 214.560 321.475 217.240 ;
        RECT 5.585 213.160 319.640 214.560 ;
        RECT 5.585 210.480 321.475 213.160 ;
        RECT 5.585 209.080 319.640 210.480 ;
        RECT 5.585 206.400 321.475 209.080 ;
        RECT 5.585 205.000 319.640 206.400 ;
        RECT 5.585 202.320 321.475 205.000 ;
        RECT 5.585 200.920 319.640 202.320 ;
        RECT 5.585 198.240 321.475 200.920 ;
        RECT 5.585 196.840 319.640 198.240 ;
        RECT 5.585 194.160 321.475 196.840 ;
        RECT 5.585 192.760 319.640 194.160 ;
        RECT 5.585 190.080 321.475 192.760 ;
        RECT 5.585 188.680 319.640 190.080 ;
        RECT 5.585 186.000 321.475 188.680 ;
        RECT 5.585 184.600 319.640 186.000 ;
        RECT 5.585 181.920 321.475 184.600 ;
        RECT 5.585 180.520 319.640 181.920 ;
        RECT 5.585 177.840 321.475 180.520 ;
        RECT 5.585 176.440 319.640 177.840 ;
        RECT 5.585 173.760 321.475 176.440 ;
        RECT 5.585 172.360 319.640 173.760 ;
        RECT 5.585 169.680 321.475 172.360 ;
        RECT 5.585 168.280 319.640 169.680 ;
        RECT 5.585 165.600 321.475 168.280 ;
        RECT 5.585 164.200 319.640 165.600 ;
        RECT 5.585 161.520 321.475 164.200 ;
        RECT 5.585 160.120 319.640 161.520 ;
        RECT 5.585 157.440 321.475 160.120 ;
        RECT 5.585 156.040 319.640 157.440 ;
        RECT 5.585 153.360 321.475 156.040 ;
        RECT 5.585 151.960 319.640 153.360 ;
        RECT 5.585 149.280 321.475 151.960 ;
        RECT 5.585 147.880 319.640 149.280 ;
        RECT 5.585 145.200 321.475 147.880 ;
        RECT 5.585 143.800 319.640 145.200 ;
        RECT 5.585 141.120 321.475 143.800 ;
        RECT 5.585 139.720 319.640 141.120 ;
        RECT 5.585 137.040 321.475 139.720 ;
        RECT 5.585 135.640 319.640 137.040 ;
        RECT 5.585 132.960 321.475 135.640 ;
        RECT 5.585 131.560 319.640 132.960 ;
        RECT 5.585 128.880 321.475 131.560 ;
        RECT 5.585 127.480 319.640 128.880 ;
        RECT 5.585 124.800 321.475 127.480 ;
        RECT 5.585 123.400 319.640 124.800 ;
        RECT 5.585 120.720 321.475 123.400 ;
        RECT 5.585 119.320 319.640 120.720 ;
        RECT 5.585 116.640 321.475 119.320 ;
        RECT 5.585 115.240 319.640 116.640 ;
        RECT 5.585 112.560 321.475 115.240 ;
        RECT 5.585 111.160 319.640 112.560 ;
        RECT 5.585 108.480 321.475 111.160 ;
        RECT 5.585 107.080 319.640 108.480 ;
        RECT 5.585 104.400 321.475 107.080 ;
        RECT 5.585 103.000 319.640 104.400 ;
        RECT 5.585 100.320 321.475 103.000 ;
        RECT 5.585 98.920 319.640 100.320 ;
        RECT 5.585 96.240 321.475 98.920 ;
        RECT 5.585 94.840 319.640 96.240 ;
        RECT 5.585 92.160 321.475 94.840 ;
        RECT 5.585 90.760 319.640 92.160 ;
        RECT 5.585 88.080 321.475 90.760 ;
        RECT 5.585 86.680 319.640 88.080 ;
        RECT 5.585 84.000 321.475 86.680 ;
        RECT 5.585 82.600 319.640 84.000 ;
        RECT 5.585 79.920 321.475 82.600 ;
        RECT 5.585 78.520 319.640 79.920 ;
        RECT 5.585 75.840 321.475 78.520 ;
        RECT 5.585 74.440 319.640 75.840 ;
        RECT 5.585 71.760 321.475 74.440 ;
        RECT 5.585 70.360 319.640 71.760 ;
        RECT 5.585 67.680 321.475 70.360 ;
        RECT 5.585 66.280 319.640 67.680 ;
        RECT 5.585 63.600 321.475 66.280 ;
        RECT 5.585 62.200 319.640 63.600 ;
        RECT 5.585 59.520 321.475 62.200 ;
        RECT 5.585 58.120 319.640 59.520 ;
        RECT 5.585 55.440 321.475 58.120 ;
        RECT 5.585 54.040 319.640 55.440 ;
        RECT 5.585 51.360 321.475 54.040 ;
        RECT 5.585 49.960 319.640 51.360 ;
        RECT 5.585 47.280 321.475 49.960 ;
        RECT 5.585 45.880 319.640 47.280 ;
        RECT 5.585 43.200 321.475 45.880 ;
        RECT 5.585 41.800 319.640 43.200 ;
        RECT 5.585 39.120 321.475 41.800 ;
        RECT 5.585 37.720 319.640 39.120 ;
        RECT 5.585 35.040 321.475 37.720 ;
        RECT 5.585 33.640 319.640 35.040 ;
        RECT 5.585 30.960 321.475 33.640 ;
        RECT 5.585 29.560 319.640 30.960 ;
        RECT 5.585 26.880 321.475 29.560 ;
        RECT 5.585 25.480 319.640 26.880 ;
        RECT 5.585 22.800 321.475 25.480 ;
        RECT 5.585 21.400 319.640 22.800 ;
        RECT 5.585 18.720 321.475 21.400 ;
        RECT 5.585 17.320 319.640 18.720 ;
        RECT 5.585 14.640 321.475 17.320 ;
        RECT 5.585 13.240 319.640 14.640 ;
        RECT 5.585 10.560 321.475 13.240 ;
        RECT 5.585 9.160 319.640 10.560 ;
        RECT 5.585 6.480 321.475 9.160 ;
        RECT 5.585 5.615 319.640 6.480 ;
      LAYER met4 ;
        RECT 10.415 11.735 20.640 296.985 ;
        RECT 23.040 11.735 97.440 296.985 ;
        RECT 99.840 11.735 174.240 296.985 ;
        RECT 176.640 11.735 251.040 296.985 ;
        RECT 253.440 11.735 310.665 296.985 ;
  END
END wb_RAxM
END LIBRARY

