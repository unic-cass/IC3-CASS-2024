magic
tech sky130A
magscale 1 2
timestamp 1731077216
<< nwell >>
rect 1066 97093 98846 97414
rect 1066 96005 98846 96571
rect 1066 94917 98846 95483
rect 1066 93829 98846 94395
rect 1066 92741 98846 93307
rect 1066 91653 98846 92219
rect 1066 90565 98846 91131
rect 1066 89477 98846 90043
rect 1066 88389 98846 88955
rect 1066 87301 98846 87867
rect 1066 86213 98846 86779
rect 1066 85125 98846 85691
rect 1066 84037 98846 84603
rect 1066 82949 98846 83515
rect 1066 81861 98846 82427
rect 1066 80773 98846 81339
rect 1066 79685 98846 80251
rect 1066 78597 98846 79163
rect 1066 77509 98846 78075
rect 1066 76421 98846 76987
rect 1066 75333 98846 75899
rect 1066 74245 98846 74811
rect 1066 73157 98846 73723
rect 1066 72069 98846 72635
rect 1066 70981 98846 71547
rect 1066 69893 98846 70459
rect 1066 68805 98846 69371
rect 1066 67717 98846 68283
rect 1066 66629 98846 67195
rect 1066 65541 98846 66107
rect 1066 64453 98846 65019
rect 1066 63365 98846 63931
rect 1066 62277 98846 62843
rect 1066 61189 98846 61755
rect 1066 60101 98846 60667
rect 1066 59013 98846 59579
rect 1066 57925 98846 58491
rect 1066 56837 98846 57403
rect 1066 55749 98846 56315
rect 1066 54661 98846 55227
rect 1066 53573 98846 54139
rect 1066 52485 98846 53051
rect 1066 51397 98846 51963
rect 1066 50309 98846 50875
rect 1066 49221 98846 49787
rect 1066 48133 98846 48699
rect 1066 47045 98846 47611
rect 1066 45957 98846 46523
rect 1066 44869 98846 45435
rect 1066 43781 98846 44347
rect 1066 42693 98846 43259
rect 1066 41605 98846 42171
rect 1066 40517 98846 41083
rect 1066 39429 98846 39995
rect 1066 38341 98846 38907
rect 1066 37253 98846 37819
rect 1066 36165 98846 36731
rect 1066 35077 98846 35643
rect 1066 33989 98846 34555
rect 1066 32901 98846 33467
rect 1066 31813 98846 32379
rect 1066 30725 98846 31291
rect 1066 29637 98846 30203
rect 1066 28549 98846 29115
rect 1066 27461 98846 28027
rect 1066 26373 98846 26939
rect 1066 25285 98846 25851
rect 1066 24197 98846 24763
rect 1066 23109 98846 23675
rect 1066 22021 98846 22587
rect 1066 20933 98846 21499
rect 1066 19845 98846 20411
rect 1066 18757 98846 19323
rect 1066 17669 98846 18235
rect 1066 16581 98846 17147
rect 1066 15493 98846 16059
rect 1066 14405 98846 14971
rect 1066 13317 98846 13883
rect 1066 12229 98846 12795
rect 1066 11141 98846 11707
rect 1066 10053 98846 10619
rect 1066 8965 98846 9531
rect 1066 7877 98846 8443
rect 1066 6789 98846 7355
rect 1066 5701 98846 6267
rect 1066 4613 98846 5179
rect 1066 3525 98846 4091
rect 1066 2437 98846 3003
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 1104 2128 98886 97424
<< metal2 >>
rect 49974 0 50030 800
<< obsm2 >>
rect 4214 856 98882 97413
rect 4214 800 49918 856
rect 50086 800 98882 856
<< metal3 >>
rect 99200 96024 100000 96144
rect 99200 91400 100000 91520
rect 99200 86776 100000 86896
rect 99200 82152 100000 82272
rect 99200 77528 100000 77648
rect 99200 72904 100000 73024
rect 99200 68280 100000 68400
rect 99200 63656 100000 63776
rect 99200 59032 100000 59152
rect 99200 54408 100000 54528
rect 99200 49784 100000 49904
rect 99200 45160 100000 45280
rect 99200 40536 100000 40656
rect 99200 35912 100000 36032
rect 99200 31288 100000 31408
rect 99200 26664 100000 26784
rect 99200 22040 100000 22160
rect 99200 17416 100000 17536
rect 99200 12792 100000 12912
rect 99200 8168 100000 8288
rect 99200 3544 100000 3664
<< obsm3 >>
rect 4210 96224 99200 97409
rect 4210 95944 99120 96224
rect 4210 91600 99200 95944
rect 4210 91320 99120 91600
rect 4210 86976 99200 91320
rect 4210 86696 99120 86976
rect 4210 82352 99200 86696
rect 4210 82072 99120 82352
rect 4210 77728 99200 82072
rect 4210 77448 99120 77728
rect 4210 73104 99200 77448
rect 4210 72824 99120 73104
rect 4210 68480 99200 72824
rect 4210 68200 99120 68480
rect 4210 63856 99200 68200
rect 4210 63576 99120 63856
rect 4210 59232 99200 63576
rect 4210 58952 99120 59232
rect 4210 54608 99200 58952
rect 4210 54328 99120 54608
rect 4210 49984 99200 54328
rect 4210 49704 99120 49984
rect 4210 45360 99200 49704
rect 4210 45080 99120 45360
rect 4210 40736 99200 45080
rect 4210 40456 99120 40736
rect 4210 36112 99200 40456
rect 4210 35832 99120 36112
rect 4210 31488 99200 35832
rect 4210 31208 99120 31488
rect 4210 26864 99200 31208
rect 4210 26584 99120 26864
rect 4210 22240 99200 26584
rect 4210 21960 99120 22240
rect 4210 17616 99200 21960
rect 4210 17336 99120 17616
rect 4210 12992 99200 17336
rect 4210 12712 99120 12992
rect 4210 8368 99200 12712
rect 4210 8088 99120 8368
rect 4210 3744 99200 8088
rect 4210 3464 99120 3744
rect 4210 2143 99200 3464
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< labels >>
rlabel metal3 s 99200 3544 100000 3664 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 99200 17416 100000 17536 6 io_in[1]
port 2 nsew signal input
rlabel metal3 s 99200 31288 100000 31408 6 io_in[2]
port 3 nsew signal input
rlabel metal3 s 99200 45160 100000 45280 6 io_in[3]
port 4 nsew signal input
rlabel metal3 s 99200 59032 100000 59152 6 io_in[4]
port 5 nsew signal input
rlabel metal3 s 99200 72904 100000 73024 6 io_in[5]
port 6 nsew signal input
rlabel metal3 s 99200 86776 100000 86896 6 io_in[6]
port 7 nsew signal input
rlabel metal3 s 99200 12792 100000 12912 6 io_oeb[0]
port 8 nsew signal output
rlabel metal3 s 99200 26664 100000 26784 6 io_oeb[1]
port 9 nsew signal output
rlabel metal3 s 99200 40536 100000 40656 6 io_oeb[2]
port 10 nsew signal output
rlabel metal3 s 99200 54408 100000 54528 6 io_oeb[3]
port 11 nsew signal output
rlabel metal3 s 99200 68280 100000 68400 6 io_oeb[4]
port 12 nsew signal output
rlabel metal3 s 99200 82152 100000 82272 6 io_oeb[5]
port 13 nsew signal output
rlabel metal3 s 99200 96024 100000 96144 6 io_oeb[6]
port 14 nsew signal output
rlabel metal3 s 99200 8168 100000 8288 6 io_out[0]
port 15 nsew signal output
rlabel metal3 s 99200 22040 100000 22160 6 io_out[1]
port 16 nsew signal output
rlabel metal3 s 99200 35912 100000 36032 6 io_out[2]
port 17 nsew signal output
rlabel metal3 s 99200 49784 100000 49904 6 io_out[3]
port 18 nsew signal output
rlabel metal3 s 99200 63656 100000 63776 6 io_out[4]
port 19 nsew signal output
rlabel metal3 s 99200 77528 100000 77648 6 io_out[5]
port 20 nsew signal output
rlabel metal3 s 99200 91400 100000 91520 6 io_out[6]
port 21 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 23 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 23 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 23 nsew ground bidirectional
rlabel metal2 s 49974 0 50030 800 6 wb_clk_i
port 24 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3452538
string GDS_FILE /media/jm/128GB_SSD/IC3-CASS-2024/openlane/user_proj_example/runs/24_11_08_11_44/results/signoff/user_proj_example.magic.gds
string GDS_START 225904
<< end >>

