* NGSPICE file created from wb_RAxM.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

.subckt wb_RAxM la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35]
+ la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40]
+ la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
+ la_data_in[47] la_data_in[4] la_data_in[5] la_data_in[6] la_data_in[7] la_data_in[8]
+ la_data_in[9] la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[3] la_data_out[4]
+ la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9] vccd2
+ vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sta_o wbs_stb_i wbs_we_i
XFILLER_0_94_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6914_ _6855_/A _7255_/B _6856_/A _6853_/Y vssd2 vssd2 vccd2 vccd2 _6914_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_89_494 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6845_ _6782_/A _6784_/B _6782_/B vssd2 vssd2 vccd2 vccd2 _6847_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__6917__B1 _6855_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_9_411 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_91_125 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6776_ _6776_/A _6776_/B _6776_/C vssd2 vssd2 vccd2 vccd2 _6776_/X sky130_fd_sc_hd__and3_1
XFILLER_0_45_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_9_466 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3988_ _3965_/A _7775_/Q _4656_/A vssd2 vssd2 vccd2 vccd2 _3988_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_91_169 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5727_ _7872_/Q _7871_/Q _5735_/B vssd2 vssd2 vccd2 vccd2 _5734_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_17_244 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_60_512 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_32_214 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_103_614 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_60_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5658_ _6019_/C _5811_/B vssd2 vssd2 vccd2 vccd2 _5658_/Y sky130_fd_sc_hd__nor2_1
X_4609_ _4609_/A _4609_/B vssd2 vssd2 vccd2 vccd2 _4610_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_60_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5589_ _5581_/A _5581_/B _5581_/C _5581_/D _5645_/B vssd2 vssd2 vccd2 vccd2 _5598_/B
+ sky130_fd_sc_hd__o41a_4
X_7328_ _7334_/C _7328_/B vssd2 vssd2 vccd2 vccd2 _7835_/D sky130_fd_sc_hd__xnor2_1
Xhold362 hold678/X vssd2 vssd2 vccd2 vccd2 _7785_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 _7752_/Q vssd2 vssd2 vccd2 vccd2 hold351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold340 _7479_/X vssd2 vssd2 vccd2 vccd2 _7719_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_472 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7259_ _7259_/A _7259_/B _7259_/C vssd2 vssd2 vccd2 vccd2 _7260_/B sky130_fd_sc_hd__and3_1
Xhold384 hold685/X vssd2 vssd2 vccd2 vccd2 _7798_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 _7683_/Q vssd2 vssd2 vccd2 vccd2 hold395/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 _7692_/Q vssd2 vssd2 vccd2 vccd2 hold373/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4459__A1 _4328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4459__B2 _4162_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4267__D _4267_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_99_225 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4564__B _4966_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_95_420 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_68_656 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_23_18 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_23_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7367__S _7383_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_82_136 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_82_103 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_36_542 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_51_512 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_23_269 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6439__A2 _7197_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4870__A1 _4966_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_442 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4960_ _4959_/B _4960_/B vssd2 vssd2 vccd2 vccd2 _4961_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_86_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_58_155 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4891_ _5164_/A _5315_/B _5105_/B _4962_/A vssd2 vssd2 vccd2 vccd2 _4891_/Y sky130_fd_sc_hd__o22ai_1
X_3911_ _3954_/C _3910_/B _3910_/C _3910_/D _4050_/B vssd2 vssd2 vccd2 vccd2 _3913_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_0_104_53 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6630_ _5819_/B _7197_/B _6627_/X vssd2 vssd2 vccd2 vccd2 _6689_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_73_125 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3842_ _7795_/Q _7796_/Q _3822_/A _3888_/B vssd2 vssd2 vccd2 vccd2 _3847_/B sky130_fd_sc_hd__o31a_2
XFILLER_0_104_97 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6561_ _6561_/A _6561_/B vssd2 vssd2 vccd2 vccd2 _6563_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_542 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_39_391 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_14_214 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5512_ _5512_/A _5512_/B vssd2 vssd2 vccd2 vccd2 _5513_/B sky130_fd_sc_hd__and2_1
X_6492_ _6855_/A _6572_/B _6415_/X _6417_/B vssd2 vssd2 vccd2 vccd2 _6502_/A sky130_fd_sc_hd__o31ai_4
XFILLER_0_89_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_42_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_112_433 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5443_ _5443_/A _5443_/B vssd2 vssd2 vccd2 vccd2 _5518_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_477 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5374_ _5431_/A _5374_/B _5468_/A _5528_/B vssd2 vssd2 vccd2 vccd2 _5417_/A sky130_fd_sc_hd__or4_1
XFILLER_0_100_628 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7113_ _7114_/A _7114_/B _7114_/C vssd2 vssd2 vccd2 vccd2 _7168_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_22_291 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4325_ _4162_/A _4519_/B _3820_/Y _4745_/A _7768_/Q vssd2 vssd2 vccd2 vccd2 _4325_/X
+ sky130_fd_sc_hd__a32o_1
X_7044_ _7197_/A _7222_/A _7222_/C _7094_/A vssd2 vssd2 vccd2 vccd2 _7046_/A sky130_fd_sc_hd__a22o_1
XANTENNA__5102__A2 _5222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4256_ _4254_/Y _4255_/X _4814_/B vssd2 vssd2 vccd2 vccd2 _4256_/X sky130_fd_sc_hd__o21a_1
X_4187_ _4187_/A _4189_/C _4189_/D vssd2 vssd2 vccd2 vccd2 _4242_/A sky130_fd_sc_hd__nand3_1
XTAP_1129 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_80 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6880__A _7037_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_77_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7877_ _7878_/CLK _7877_/D _7636_/Y vssd2 vssd2 vccd2 vccd2 _7877_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_37_306 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6366__A1 _6668_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6828_ _6829_/A _6829_/B vssd2 vssd2 vccd2 vccd2 _6828_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_49_188 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_37_328 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_107_205 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_92_456 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_18_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_107_249 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6759_ _6693_/A _6693_/B _6691_/Y vssd2 vssd2 vccd2 vccd2 _6763_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_92_489 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_60_331 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_20_206 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_444 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_20_239 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold170 _7433_/X vssd2 vssd2 vccd2 vccd2 _7434_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _7361_/X vssd2 vssd2 vccd2 vccd2 _7362_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _7355_/X vssd2 vssd2 vccd2 vccd2 _7356_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1630 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_95_261 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_83_412 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4741__C _4965_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_158 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_50_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_83_489 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_24_567 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_24_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5090_ _5091_/A _5091_/B _5089_/Y vssd2 vssd2 vccd2 vccd2 _5090_/X sky130_fd_sc_hd__o21ba_1
X_4110_ _7767_/Q _4458_/D vssd2 vssd2 vccd2 vccd2 _4110_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4041_ _4454_/A _4122_/D _4066_/C _4066_/D vssd2 vssd2 vccd2 vccd2 _4041_/X sky130_fd_sc_hd__and4_1
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_420 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7800_ _7800_/CLK _7800_/D _7559_/Y vssd2 vssd2 vccd2 vccd2 _7800_/Q sky130_fd_sc_hd__dfrtp_4
X_5992_ _6510_/A _5992_/B _5992_/C vssd2 vssd2 vccd2 vccd2 _5992_/X sky130_fd_sc_hd__and3_1
X_4943_ _4943_/A _4943_/B vssd2 vssd2 vccd2 vccd2 _4946_/A sky130_fd_sc_hd__xnor2_1
X_7731_ _7776_/CLK _7731_/D _7490_/Y vssd2 vssd2 vccd2 vccd2 _7731_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7662_ _7806_/CLK _7662_/D vssd2 vssd2 vccd2 vccd2 _7662_/Q sky130_fd_sc_hd__dfxtp_1
X_6613_ _6613_/A _6613_/B vssd2 vssd2 vccd2 vccd2 _6765_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__6205__A _6634_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4874_ _4874_/A _4874_/B vssd2 vssd2 vccd2 vccd2 _4876_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_467 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7593_ _7597_/A vssd2 vssd2 vccd2 vccd2 _7593_/Y sky130_fd_sc_hd__inv_2
X_3825_ _7805_/Q _3825_/B vssd2 vssd2 vccd2 vccd2 _5458_/A sky130_fd_sc_hd__xnor2_4
X_6544_ _5778_/X _5786_/Y _7253_/B _5736_/X vssd2 vssd2 vccd2 vccd2 _6547_/A sky130_fd_sc_hd__a211o_1
XFILLER_0_61_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_383 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6475_ _6550_/A _6636_/A _7253_/A _7253_/B vssd2 vssd2 vccd2 vccd2 _6542_/A sky130_fd_sc_hd__or4_2
XFILLER_0_42_342 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_15_556 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_30_504 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_40_93 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5426_ _5427_/B _5427_/A vssd2 vssd2 vccd2 vccd2 _5480_/A sky130_fd_sc_hd__and2b_1
XANTENNA__4379__B _5220_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5357_ _5357_/A _5357_/B _5357_/C _5257_/A vssd2 vssd2 vccd2 vccd2 _5454_/B sky130_fd_sc_hd__or4b_2
X_5288_ _5289_/A _5289_/B vssd2 vssd2 vccd2 vccd2 _5288_/Y sky130_fd_sc_hd__nand2b_1
X_4308_ _4308_/A _4308_/B vssd2 vssd2 vccd2 vccd2 _4309_/B sky130_fd_sc_hd__nand2_1
X_7027_ _6762_/A _6836_/Y _6838_/B _7025_/C _7025_/D vssd2 vssd2 vccd2 vccd2 _7029_/A
+ sky130_fd_sc_hd__a2111o_1
X_4239_ _4239_/A _4239_/B vssd2 vssd2 vccd2 vccd2 _4243_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_90 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_108_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_53_607 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_37_136 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_92_253 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_80_415 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_404 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_37_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_80_459 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_20_19 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_45_191 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_21_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5314__A2 _5498_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_29_28 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_88_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_88_537 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_15 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1460 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_581 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1493 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_220 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_83_264 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_114_517 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4590_ _4662_/B _5042_/B _5222_/A _4962_/A vssd2 vssd2 vccd2 vccd2 _4590_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_43_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_24_331 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_397 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6260_ _6261_/A _6261_/B _6261_/C vssd2 vssd2 vccd2 vccd2 _6381_/A sky130_fd_sc_hd__o21a_2
X_5211_ _5211_/A _5211_/B vssd2 vssd2 vccd2 vccd2 _5213_/A sky130_fd_sc_hd__nand2_1
X_6191_ _6398_/A _6253_/B _6191_/C _6191_/D vssd2 vssd2 vccd2 vccd2 _6191_/X sky130_fd_sc_hd__and4_1
X_5142_ _5207_/A _5431_/A _5142_/C _5498_/A vssd2 vssd2 vccd2 vccd2 _5201_/A sky130_fd_sc_hd__or4_2
XFILLER_0_19_50 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5073_ _5042_/A _5431_/B _5192_/A _5072_/Y vssd2 vssd2 vccd2 vccd2 _5119_/A sky130_fd_sc_hd__o22ai_4
XFILLER_0_79_515 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4024_ _4893_/A _4315_/B _4427_/A vssd2 vssd2 vccd2 vccd2 _4025_/C sky130_fd_sc_hd__and3_1
XANTENNA__6580__D _7224_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5975_ _6158_/A _5791_/X _5825_/X _6074_/A vssd2 vssd2 vccd2 vccd2 _5975_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_47_456 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_47_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4926_ _4926_/A _4997_/B vssd2 vssd2 vccd2 vccd2 _7742_/D sky130_fd_sc_hd__xnor2_1
X_7714_ _7771_/CLK _7714_/D vssd2 vssd2 vccd2 vccd2 _7714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_125 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4857_ _4598_/A _5431_/B _4855_/Y vssd2 vssd2 vccd2 vccd2 _4916_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_51_70 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7645_ _7645_/A vssd2 vssd2 vccd2 vccd2 _7645_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_670 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7576_ _7590_/A vssd2 vssd2 vccd2 vccd2 _7576_/Y sky130_fd_sc_hd__inv_2
X_3808_ _7799_/Q _7800_/Q _3822_/A _3822_/B _3888_/B vssd2 vssd2 vccd2 vccd2 _3831_/B
+ sky130_fd_sc_hd__o41a_4
X_6527_ _6527_/A _6527_/B vssd2 vssd2 vccd2 vccd2 _6528_/B sky130_fd_sc_hd__xnor2_2
X_4788_ _4789_/A _4789_/B vssd2 vssd2 vccd2 vccd2 _4788_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__6589__B _7313_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_43_651 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_70_481 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_113_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6458_ _6615_/A vssd2 vssd2 vccd2 vccd2 _6458_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_100_233 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6389_ _6389_/A _6389_/B vssd2 vssd2 vccd2 vccd2 _6390_/C sky130_fd_sc_hd__or2_1
X_5409_ _5475_/A _5475_/B vssd2 vssd2 vccd2 vccd2 _5476_/A sky130_fd_sc_hd__or2_1
XFILLER_0_100_277 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5014__A _5210_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7221__A2 _7253_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_78_570 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_108_333 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_38_489 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_108_377 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_93_595 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7375__S _7383_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_25_117 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_108_399 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_104_583 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_104_594 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_507 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_56_59 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_88_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__7460__A2 _7454_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_72_47 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_88_378 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_76_529 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_69_592 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_8_328 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5760_ _5760_/A _5760_/B _5760_/C _5760_/D vssd2 vssd2 vccd2 vccd2 _5760_/X sky130_fd_sc_hd__or4_1
XANTENNA__6971__A1 _6571_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1290 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4711_ _4711_/A _5042_/B _4782_/B _5099_/A vssd2 vssd2 vccd2 vccd2 _4712_/B sky130_fd_sc_hd__or4_1
X_5691_ _5691_/A _5691_/B vssd2 vssd2 vccd2 vccd2 _6281_/B sky130_fd_sc_hd__and2_4
XFILLER_0_112_53 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4642_ _4643_/B _4643_/A vssd2 vssd2 vccd2 vccd2 _4642_/X sky130_fd_sc_hd__and2b_1
X_7430_ _7436_/A _7430_/B vssd2 vssd2 vccd2 vccd2 _7683_/D sky130_fd_sc_hd__and2_1
XFILLER_0_112_97 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4573_ _4573_/A _4573_/B vssd2 vssd2 vccd2 vccd2 _4610_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_52_470 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4734__B1 _5374_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7361_ hold180/X _7651_/Q _7383_/S vssd2 vssd2 vccd2 vccd2 _7361_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_673 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_31_109 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_97_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6312_ _6181_/Y _6308_/B _6311_/C _6184_/X vssd2 vssd2 vccd2 vccd2 _6313_/C sky130_fd_sc_hd__o22a_1
X_7292_ _7253_/B _7253_/D _6670_/Y _7253_/A vssd2 vssd2 vccd2 vccd2 _7292_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_12_323 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_24_183 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6243_ _6177_/A _6177_/B _6175_/X vssd2 vssd2 vccd2 vccd2 _6245_/B sky130_fd_sc_hd__a21oi_2
X_6174_ _6115_/A _6115_/C _6115_/B vssd2 vssd2 vccd2 vccd2 _6176_/B sky130_fd_sc_hd__o21ba_1
X_5125_ _5126_/A _5126_/B vssd2 vssd2 vccd2 vccd2 _5125_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_98_109 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5056_ _5056_/A _5056_/B vssd2 vssd2 vccd2 vccd2 _5059_/A sky130_fd_sc_hd__xnor2_4
X_4007_ _4149_/B _4149_/C vssd2 vssd2 vccd2 vccd2 _4075_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_67_529 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_94_359 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_94_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5958_ _5958_/A _5958_/B _5958_/C vssd2 vssd2 vccd2 vccd2 _5960_/A sky130_fd_sc_hd__and3_1
XFILLER_0_62_91 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_47_220 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4909_ _4826_/A _4826_/B _4824_/Y vssd2 vssd2 vccd2 vccd2 _4911_/B sky130_fd_sc_hd__a21bo_2
XFILLER_0_47_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_404 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_75_584 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_62_201 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5889_ _5883_/A _5875_/X _5883_/C _5888_/X _6424_/A vssd2 vssd2 vccd2 vccd2 _5890_/B
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_90_554 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7628_ _7629_/A vssd2 vssd2 vccd2 vccd2 _7628_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_105_369 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_62_278 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_43_481 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7559_ _7563_/A vssd2 vssd2 vccd2 vccd2 _7559_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5009__A _5168_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_113_391 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6478__B1 _6404_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_31_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7224__A _7224_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4848__A _4849_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold30 hold30/A vssd2 vssd2 vccd2 vccd2 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd2 vssd2 vccd2 vccd2 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd2 vssd2 vccd2 vccd2 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd2 vssd2 vccd2 vccd2 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd2 vssd2 vccd2 vccd2 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4341__A_N _5042_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold96 hold96/A vssd2 vssd2 vccd2 vccd2 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd2 vssd2 vccd2 vccd2 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5756__A2 _5781_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_66_573 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_38_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_38_264 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_108_141 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_26_448 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_81_543 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_14_wb_clk_i clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7787_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_317 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA_5 wbs_adr_i[11] vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5861__B _6707_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_1_537 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_315 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5141__B1 _5498_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_348 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4495__A2 _4711_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6973__A _6973_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_359 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4493__A _4598_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5995__A2 _5993_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6930_ _6930_/A _6930_/B vssd2 vssd2 vccd2 vccd2 _6932_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_16_40 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_76_304 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6861_ _7047_/A _7145_/A vssd2 vssd2 vccd2 vccd2 _6862_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_88_197 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6792_ _6793_/A _6793_/B vssd2 vssd2 vccd2 vccd2 _6792_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_9_604 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5812_ _6093_/A _6424_/A _5812_/C _5812_/D vssd2 vssd2 vccd2 vccd2 _5812_/X sky130_fd_sc_hd__and4_1
X_5743_ _6587_/A _6510_/B _6670_/B vssd2 vssd2 vccd2 vccd2 _5744_/B sky130_fd_sc_hd__or3_4
XFILLER_0_29_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_91_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_84_392 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4940__B _5210_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_57_584 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_17_415 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_32_61 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6213__A _6855_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5674_ _5674_/A _5674_/B _5674_/C _5674_/D vssd2 vssd2 vccd2 vccd2 _5674_/X sky130_fd_sc_hd__or4_2
X_4625_ _4570_/A _4570_/B _4568_/Y vssd2 vssd2 vccd2 vccd2 _4643_/A sky130_fd_sc_hd__a21o_1
X_7413_ _7452_/A _7413_/B vssd2 vssd2 vccd2 vccd2 _7675_/D sky130_fd_sc_hd__and2_1
XFILLER_0_32_429 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold511 hold40/X vssd2 vssd2 vccd2 vccd2 _7854_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7344_ _7344_/A _7344_/B _7344_/C _7344_/D vssd2 vssd2 vccd2 vccd2 _7345_/D sky130_fd_sc_hd__or4_1
X_4556_ _4556_/A _4556_/B vssd2 vssd2 vccd2 vccd2 _4557_/B sky130_fd_sc_hd__or2_1
Xhold500 la_data_in[27] vssd2 vssd2 vccd2 vccd2 hold47/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 la_data_in[45] vssd2 vssd2 vccd2 vccd2 hold69/A sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap241 _4326_/D vssd2 vssd2 vccd2 vccd2 _4268_/D sky130_fd_sc_hd__buf_2
XFILLER_0_12_164 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold522 input11/X vssd2 vssd2 vccd2 vccd2 hold76/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3930__A1 _7762_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold533 hold57/X vssd2 vssd2 vccd2 vccd2 input18/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_440 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7275_ _7275_/A _7275_/B vssd2 vssd2 vccd2 vccd2 _7277_/B sky130_fd_sc_hd__or2_1
Xhold555 hold68/X vssd2 vssd2 vccd2 vccd2 _7851_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4487_ _4452_/A _4452_/B _4450_/Y vssd2 vssd2 vccd2 vccd2 _4504_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_12_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold577 hold81/X vssd2 vssd2 vccd2 vccd2 input45/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 la_data_in[5] vssd2 vssd2 vccd2 vccd2 hold87/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 input14/X vssd2 vssd2 vccd2 vccd2 hold66/A sky130_fd_sc_hd__dlygate4sd3_1
X_6226_ _6590_/A _7197_/A vssd2 vssd2 vccd2 vccd2 _6228_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4387__B _4965_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold599 hold92/X vssd2 vssd2 vccd2 vccd2 _7874_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_871 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6157_/A _6510_/B vssd2 vssd2 vccd2 vccd2 _6157_/X sky130_fd_sc_hd__and2_1
X_5108_ _5048_/A _5048_/B _5046_/X vssd2 vssd2 vccd2 vccd2 _5110_/B sky130_fd_sc_hd__o21a_2
XTAP_893 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6088_ _6634_/B _6664_/A _5948_/X _5931_/C vssd2 vssd2 vccd2 vccd2 _6090_/A sky130_fd_sc_hd__a22o_1
X_5039_ _5164_/A _5468_/A _5550_/B _4962_/A vssd2 vssd2 vccd2 vccd2 _5048_/A sky130_fd_sc_hd__o22a_2
XANTENNA__5011__B _5550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_67_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_82_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6935__A1 _6039_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7219__A _7336_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_94_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_63_510 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_212 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_656 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_105_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_90_373 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_63_587 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_50_237 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4174__A1 _4044_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5457__A2_N _5498_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_31_462 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4463__D _5099_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XPHY_170 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_54_521 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_192 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_181 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6033__A _6092_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_54_543 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4410_ _4291_/A _4291_/B _4351_/B _4352_/B _4352_/A vssd2 vssd2 vccd2 vccd2 _4412_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_112_637 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_111_125 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5390_ _5390_/A _5390_/B vssd2 vssd2 vccd2 vccd2 _5392_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_111_169 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_78_79 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4341_ _5042_/A _5030_/B _5030_/A vssd2 vssd2 vccd2 vccd2 _4345_/A sky130_fd_sc_hd__and3b_2
XFILLER_0_1_367 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7060_ _7060_/A _7060_/B vssd2 vssd2 vccd2 vccd2 _7062_/B sky130_fd_sc_hd__xnor2_1
X_4272_ _4810_/A _5042_/B vssd2 vssd2 vccd2 vccd2 _4277_/A sky130_fd_sc_hd__nor2_2
X_6011_ _6011_/A _6068_/B vssd2 vssd2 vccd2 vccd2 _7812_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_27_72 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_89_462 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6913_ _6775_/X _6901_/B _6899_/X vssd2 vssd2 vccd2 vccd2 _6967_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_76_123 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_49_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_49_326 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6844_ _6798_/A _6798_/B _6796_/X vssd2 vssd2 vccd2 vccd2 _6847_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_64_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6917__B2 _7291_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6775_ _6776_/A _6776_/B _6776_/C vssd2 vssd2 vccd2 vccd2 _6775_/X sky130_fd_sc_hd__a21o_1
X_3987_ _4033_/C _4125_/C _4057_/C vssd2 vssd2 vccd2 vccd2 _3987_/X sky130_fd_sc_hd__and3_1
XFILLER_0_91_137 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_72_340 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5726_ _6100_/D _6587_/B _5938_/C _5898_/C vssd2 vssd2 vccd2 vccd2 _5992_/C sky130_fd_sc_hd__and4_2
Xwb_RAxM_294 vssd2 vssd2 vccd2 vccd2 wb_RAxM_294/HI wbs_sta_o sky130_fd_sc_hd__conb_1
XFILLER_0_5_673 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5782__A _6282_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5657_ _5828_/B _5828_/C _6191_/D _5630_/B _6075_/C vssd2 vssd2 vccd2 vccd2 _5921_/D
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_0_103_659 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4608_ _4609_/A _4609_/B vssd2 vssd2 vccd2 vccd2 _4608_/Y sky130_fd_sc_hd__nor2_1
X_5588_ _5586_/B _5584_/Y _5587_/X vssd2 vssd2 vccd2 vccd2 _5588_/Y sky130_fd_sc_hd__o21ai_4
X_7327_ _7335_/A _7335_/B _6069_/A vssd2 vssd2 vccd2 vccd2 _7328_/B sky130_fd_sc_hd__o21a_1
XANTENNA__4398__A _5029_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4539_ _4539_/A _4539_/B vssd2 vssd2 vccd2 vccd2 _4542_/A sky130_fd_sc_hd__xor2_2
Xhold352 _7480_/X vssd2 vssd2 vccd2 vccd2 _7720_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 _7749_/Q vssd2 vssd2 vccd2 vccd2 hold341/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold330 _7471_/X vssd2 vssd2 vccd2 vccd2 _7711_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_484 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_40_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7258_ _7259_/A _7259_/B _7259_/C vssd2 vssd2 vccd2 vccd2 _7289_/A sky130_fd_sc_hd__a21oi_1
Xhold385 _7654_/Q vssd2 vssd2 vccd2 vccd2 hold385/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 hold679/X vssd2 vssd2 vccd2 vccd2 _7763_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 hold688/X vssd2 vssd2 vccd2 vccd2 _7778_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 _7660_/Q vssd2 vssd2 vccd2 vccd2 hold396/X sky130_fd_sc_hd__dlygate4sd3_1
X_6209_ _6210_/A _6210_/B vssd2 vssd2 vccd2 vccd2 _6261_/A sky130_fd_sc_hd__and2_1
X_7189_ _7232_/B _7189_/B vssd2 vssd2 vccd2 vccd2 _7189_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5408__A1 _5366_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_690 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_237 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4564__C _4711_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_95_432 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_68_635 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_67_101 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4861__A _5042_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_82_115 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_36_554 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_63_351 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6788__A _6989_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_51_557 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_51_535 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7383__S _7383_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5895__B2 _7845_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_31_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_64_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6028__A _6812_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4870__A2 _5276_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6072__A1 _6282_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6072__B2 _7849_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_86_454 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_80_47 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4890_ _4949_/B _4890_/B vssd2 vssd2 vccd2 vccd2 _4908_/A sky130_fd_sc_hd__nor2_2
X_3910_ _3954_/C _3910_/B _3910_/C _3910_/D vssd2 vssd2 vccd2 vccd2 _3927_/B sky130_fd_sc_hd__or4_1
XFILLER_0_86_498 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3841_ _4458_/C _4141_/C vssd2 vssd2 vccd2 vccd2 _4082_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_104_65 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6560_ _6561_/B _6561_/A vssd2 vssd2 vccd2 vccd2 _6631_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_13_52 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5511_ _5512_/A _5512_/B vssd2 vssd2 vccd2 vccd2 _5541_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_112_401 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6491_ _6491_/A _6491_/B vssd2 vssd2 vccd2 vccd2 _6528_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_557 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_14_248 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5442_ _5443_/B _5443_/A vssd2 vssd2 vccd2 vccd2 _5488_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_112_445 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5373_ _5374_/B _5468_/A _5528_/B _5222_/A vssd2 vssd2 vccd2 vccd2 _5373_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_0_112_489 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7088__B1 _6669_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7112_ _7048_/A _7048_/B _7046_/B vssd2 vssd2 vccd2 vccd2 _7114_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__4011__A _7767_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4324_ _4413_/A _4324_/B vssd2 vssd2 vccd2 vccd2 _4352_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_10_454 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_10_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7043_ _6999_/A _6999_/B _7000_/Y vssd2 vssd2 vccd2 vccd2 _7062_/A sky130_fd_sc_hd__a21bo_1
X_4255_ _7767_/Q _4707_/A _4063_/X _7769_/Q vssd2 vssd2 vccd2 vccd2 _4255_/X sky130_fd_sc_hd__a22o_1
X_4186_ _4186_/A _4186_/B vssd2 vssd2 vccd2 vccd2 _4189_/D sky130_fd_sc_hd__xor2_1
XANTENNA_fanout272_A _7772_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_89_281 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1108 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6880__B _7237_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7876_ _7878_/CLK _7876_/D _7635_/Y vssd2 vssd2 vccd2 vccd2 _7876_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6366__A2 _7094_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6827_ _6750_/A _6750_/B _6748_/Y vssd2 vssd2 vccd2 vccd2 _6829_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_107_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5574__B1 _5548_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4377__A1 _4656_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6758_ _6758_/A _6758_/B vssd2 vssd2 vccd2 vccd2 _6763_/A sky130_fd_sc_hd__xnor2_2
X_6689_ _6689_/A _6689_/B vssd2 vssd2 vccd2 vccd2 _6692_/A sky130_fd_sc_hd__xnor2_2
X_5709_ _7877_/Q _5694_/A _5694_/B _5735_/B vssd2 vssd2 vccd2 vccd2 _5710_/B sky130_fd_sc_hd__o31a_2
XFILLER_0_103_423 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__6401__A _6550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_60_387 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5877__A1 _6283_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold171 wbs_dat_i[5] vssd2 vssd2 vccd2 vccd2 input94/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 hold358/X vssd2 vssd2 vccd2 vccd2 _7775_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 hold377/X vssd2 vssd2 vccd2 vccd2 _7765_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 wbs_dat_i[13] vssd2 vssd2 vccd2 vccd2 input87/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_19 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4856__A _4893_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_34_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XTAP_1631 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_465 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_68_443 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4591__A _4962_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_95_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4741__D _5406_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5565__B1 _5548_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_3_418 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_51_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__7407__A _7452_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6030__B _6738_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_75_69 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4040_ _7762_/Q _4019_/Y _4160_/B _7766_/Q _4039_/X vssd2 vssd2 vccd2 vccd2 _4040_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_59_432 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_59_410 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5991_ _5850_/B _5987_/X _5988_/X _5990_/X vssd2 vssd2 vccd2 vccd2 _5991_/X sky130_fd_sc_hd__a211o_2
XFILLER_0_86_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4942_ _5207_/A _5366_/A vssd2 vssd2 vccd2 vccd2 _4943_/B sky130_fd_sc_hd__nor2_1
X_7730_ _7739_/CLK _7730_/D _7489_/Y vssd2 vssd2 vccd2 vccd2 _7730_/Q sky130_fd_sc_hd__dfrtp_1
X_7661_ _7806_/CLK _7661_/D vssd2 vssd2 vccd2 vccd2 _7661_/Q sky130_fd_sc_hd__dfxtp_1
X_6612_ _6613_/A _6613_/B vssd2 vssd2 vccd2 vccd2 _6612_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6205__B _6571_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4873_ _4873_/A _4873_/B vssd2 vssd2 vccd2 vccd2 _4874_/B sky130_fd_sc_hd__nand2_2
X_7592_ _7597_/A vssd2 vssd2 vccd2 vccd2 _7592_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3824_ _7805_/Q _3825_/B vssd2 vssd2 vccd2 vccd2 _3824_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_104_209 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6543_ _6502_/A _6501_/B _6499_/X vssd2 vssd2 vccd2 vccd2 _6564_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_15_535 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_40_61 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6474_ _6474_/A _6474_/B vssd2 vssd2 vccd2 vccd2 _7253_/B sky130_fd_sc_hd__nand2_8
XFILLER_0_42_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__3845__A _4267_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5859__B2 _7847_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5859__A1 _6158_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5425_ _5412_/B _5380_/B _5382_/B _5382_/A vssd2 vssd2 vccd2 vccd2 _5427_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_112_253 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_100_426 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_64_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_23_590 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_100_448 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5356_ _5445_/A _5356_/B vssd2 vssd2 vccd2 vccd2 _5454_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_10_262 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5287_ _5287_/A _5287_/B vssd2 vssd2 vccd2 vccd2 _5289_/B sky130_fd_sc_hd__xnor2_2
X_4307_ _4308_/A _4307_/B vssd2 vssd2 vccd2 vccd2 _7733_/D sky130_fd_sc_hd__xnor2_1
X_7026_ _6767_/A _6767_/B _6767_/C _7025_/X vssd2 vssd2 vccd2 vccd2 _7031_/B sky130_fd_sc_hd__a31o_1
XANTENNA__7481__B1 _7483_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6284__A1 _6093_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4238_ _4181_/A _4181_/B _4179_/Y vssd2 vssd2 vccd2 vccd2 _4239_/B sky130_fd_sc_hd__a21o_1
X_4169_ _7764_/Q _4815_/B _4032_/C _7766_/Q _4168_/X vssd2 vssd2 vccd2 vccd2 _4169_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6992__C1 _7143_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_92_221 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_65_457 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7859_ _7886_/CLK _7859_/D _7618_/Y vssd2 vssd2 vccd2 vccd2 _7859_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_37_126 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_37_148 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_108_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_92_265 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_45_181 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_33_321 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_354 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5970__A _7336_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_60_184 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7472__B1 _7483_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1450 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5210__A _5210_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1483 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1494 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_276 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_56_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_71_449 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_114_529 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_101_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_12_527 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6976__A _7037_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5210_ _5210_/A _5210_/B _5528_/A _5498_/D vssd2 vssd2 vccd2 vccd2 _5211_/B sky130_fd_sc_hd__or4_1
XANTENNA__5880__A _7847_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6190_ _7336_/A _6316_/A vssd2 vssd2 vccd2 vccd2 _6250_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4496__A _4704_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5141_ _5431_/A _5142_/C _5498_/A _5099_/A vssd2 vssd2 vccd2 vccd2 _5143_/A sky130_fd_sc_hd__o22ai_1
X_5072_ _5072_/A _5072_/B _5072_/C vssd2 vssd2 vccd2 vccd2 _5072_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__7463__B1 _7485_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4023_ _4315_/B _4214_/B _4070_/D vssd2 vssd2 vccd2 vccd2 _4251_/B sky130_fd_sc_hd__and3_1
XFILLER_0_79_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7600__A _7627_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_240 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__5758__C _7846_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_35_72 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5974_ _5974_/A _5974_/B vssd2 vssd2 vccd2 vccd2 _5985_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__4662__C _5099_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7713_ _7771_/CLK _7713_/D vssd2 vssd2 vccd2 vccd2 _7713_/Q sky130_fd_sc_hd__dfxtp_1
X_4925_ _4925_/A _4925_/B vssd2 vssd2 vccd2 vccd2 _4997_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_47_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7644_ _7645_/A vssd2 vssd2 vccd2 vccd2 _7644_/Y sky130_fd_sc_hd__inv_2
X_4856_ _4893_/A _4856_/B vssd2 vssd2 vccd2 vccd2 _5431_/B sky130_fd_sc_hd__nand2_8
X_7575_ _7590_/A vssd2 vssd2 vccd2 vccd2 _7575_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_51_93 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_51_82 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_3807_ _7795_/Q _7796_/Q _7797_/Q _7798_/Q vssd2 vssd2 vccd2 vccd2 _3822_/B sky130_fd_sc_hd__or4_4
XFILLER_0_105_529 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6526_ _6527_/B _6527_/A vssd2 vssd2 vccd2 vccd2 _6526_/Y sky130_fd_sc_hd__nand2b_1
X_4787_ _4787_/A _4787_/B vssd2 vssd2 vccd2 vccd2 _4789_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_55_490 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7047__A _7047_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_15_343 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_15_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6457_ _6457_/A _6457_/B vssd2 vssd2 vccd2 vccd2 _6615_/A sky130_fd_sc_hd__xor2_2
XANTENNA__5790__A _6157_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6388_ _6387_/A _6387_/B _6387_/C vssd2 vssd2 vccd2 vccd2 _6389_/B sky130_fd_sc_hd__a21oi_1
X_5408_ _5366_/A _5550_/B _5407_/Y vssd2 vssd2 vccd2 vccd2 _5475_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_100_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5339_ _5339_/A _5339_/B vssd2 vssd2 vccd2 vccd2 _5344_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_289 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5014__B _5210_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7009_ _7010_/A _7010_/B _7008_/X vssd2 vssd2 vccd2 vccd2 _7077_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_97_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_78_582 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5030__A _5030_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_108_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_31_19 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_108_345 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_65_287 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_53_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_108_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4743__A1 _4656_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_18_181 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4743__B2 _4809_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_21_379 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_508 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4747__C _5528_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_56_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5205__A _5328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_56_49 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__6036__A _7847_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6971__A2 _7222_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1291 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_574 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4710_ _5042_/B _4782_/B _5099_/A _4711_/A vssd2 vssd2 vccd2 vccd2 _4712_/A sky130_fd_sc_hd__o22ai_1
XFILLER_0_56_265 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5875__A _7844_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5690_ _7882_/Q _5690_/B _5690_/C vssd2 vssd2 vccd2 vccd2 _5691_/B sky130_fd_sc_hd__or3_4
XFILLER_0_29_479 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4641_ _4641_/A _4641_/B vssd2 vssd2 vccd2 vccd2 _4643_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_287 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_112_65 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_114_337 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4572_ _4572_/A _4572_/B vssd2 vssd2 vccd2 vccd2 _4573_/B sky130_fd_sc_hd__xnor2_2
X_7360_ _7436_/A _7360_/B vssd2 vssd2 vccd2 vccd2 _7650_/D sky130_fd_sc_hd__and2_1
X_6311_ _6311_/A _6311_/B _6311_/C _6186_/B vssd2 vssd2 vccd2 vccd2 _6313_/B sky130_fd_sc_hd__or4b_2
X_7291_ _7291_/A _7291_/B vssd2 vssd2 vccd2 vccd2 _7297_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4003__B _5458_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6242_ _6242_/A _6242_/B vssd2 vssd2 vccd2 vccd2 _6245_/A sky130_fd_sc_hd__xnor2_2
X_6173_ _6173_/A _6173_/B vssd2 vssd2 vccd2 vccd2 _6176_/A sky130_fd_sc_hd__xor2_2
X_5124_ _5064_/A _5064_/B _5062_/Y vssd2 vssd2 vccd2 vccd2 _5126_/B sky130_fd_sc_hd__a21oi_4
X_5055_ _5055_/A _5055_/B vssd2 vssd2 vccd2 vccd2 _5056_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__4954__A _5030_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_27_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4006_ _4656_/C _4006_/B _4006_/C vssd2 vssd2 vccd2 vccd2 _4149_/C sky130_fd_sc_hd__or3_1
XFILLER_0_67_508 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_87_390 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5957_ _5956_/A _5956_/B _5956_/C vssd2 vssd2 vccd2 vccd2 _5958_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_232 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4908_ _4908_/A _4908_/B vssd2 vssd2 vccd2 vccd2 _4911_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__5785__A _6152_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_62_224 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5888_ _7843_/Q _5588_/Y _5873_/X vssd2 vssd2 vccd2 vccd2 _5888_/X sky130_fd_sc_hd__a21o_1
X_7627_ _7627_/A vssd2 vssd2 vccd2 vccd2 _7627_/Y sky130_fd_sc_hd__inv_2
X_4839_ _4839_/A _4839_/B vssd2 vssd2 vccd2 vccd2 _4841_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_337 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_62_268 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7558_ _7561_/A vssd2 vssd2 vccd2 vccd2 _7558_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5009__B _5207_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6509_ _5816_/A _5816_/B _7291_/A vssd2 vssd2 vccd2 vccd2 _6515_/A sky130_fd_sc_hd__a21oi_2
X_7489_ _7524_/A vssd2 vssd2 vccd2 vccd2 _7489_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_101_532 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6478__A1 _5948_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6478__B2 _6634_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5951__C _6783_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_30_165 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__7224__B _7255_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_101_576 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold31 hold31/A vssd2 vssd2 vccd2 vccd2 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A vssd2 vssd2 vccd2 vccd2 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd2 vssd2 vccd2 vccd2 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd2 vssd2 vccd2 vccd2 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd2 vssd2 vccd2 vccd2 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_611 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold97 wbs_adr_i[1] vssd2 vssd2 vccd2 vccd2 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd2 vssd2 vccd2 vccd2 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd2 vssd2 vccd2 vccd2 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4661__B1 _5315_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_58_519 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_109_665 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_93_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_81_522 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_109_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_108_153 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_108_197 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_22_611 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA_6 wbs_dat_i[8] vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_21_110 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_111_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__7415__A _7450_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_67_48 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_305 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5141__B2 _5099_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5141__A1 _5431_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_349 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6973__B _6973_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_83_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4493__B _5142_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_16_52 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_49_519 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6860_ _6860_/A _6860_/B vssd2 vssd2 vccd2 vccd2 _6862_/A sky130_fd_sc_hd__xnor2_1
X_6791_ _6939_/A _7181_/A _6714_/A _6711_/X vssd2 vssd2 vccd2 vccd2 _6793_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_57_530 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_29_221 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5811_ _6019_/C _5811_/B _5811_/C _5878_/B vssd2 vssd2 vccd2 vccd2 _5812_/D sky130_fd_sc_hd__nor4_1
X_5742_ _6283_/B _6094_/B _6102_/C _5742_/D vssd2 vssd2 vccd2 vccd2 _5936_/B sky130_fd_sc_hd__and4bb_2
XFILLER_0_84_371 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4940__C _5222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_57_596 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_17_427 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__6213__B _6581_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_72_566 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_72_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_17_449 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5673_ _5663_/X _5667_/X _5672_/X _5631_/X vssd2 vssd2 vccd2 vccd2 _5674_/D sky130_fd_sc_hd__a22o_1
X_4624_ _4573_/A _4573_/B _4571_/Y vssd2 vssd2 vccd2 vccd2 _4681_/A sky130_fd_sc_hd__a21bo_1
X_7412_ hold158/X _7787_/D _7418_/S vssd2 vssd2 vccd2 vccd2 _7412_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_102_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_52_290 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7343_ _7343_/A _7343_/B _7343_/C _7343_/D vssd2 vssd2 vccd2 vccd2 _7345_/C sky130_fd_sc_hd__or4_1
X_4555_ _4556_/A _4555_/B vssd2 vssd2 vccd2 vccd2 _7737_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_644 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold501 hold47/X vssd2 vssd2 vccd2 vccd2 input20/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7325__A _7334_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold545 hold69/X vssd2 vssd2 vccd2 vccd2 input40/A sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap242 _3982_/B vssd2 vssd2 vccd2 vccd2 _4856_/B sky130_fd_sc_hd__buf_4
Xhold523 hold76/X vssd2 vssd2 vccd2 vccd2 _7858_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap231 _5812_/D vssd2 vssd2 vccd2 vccd2 _5834_/B sky130_fd_sc_hd__buf_1
Xhold534 input18/X vssd2 vssd2 vccd2 vccd2 hold58/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 la_data_in[26] vssd2 vssd2 vccd2 vccd2 hold45/A sky130_fd_sc_hd__dlygate4sd3_1
X_7274_ _7303_/B _7274_/B vssd2 vssd2 vccd2 vccd2 _7277_/A sky130_fd_sc_hd__nor2_1
X_4486_ _4441_/A _4441_/B _4439_/X vssd2 vssd2 vccd2 vccd2 _4543_/A sky130_fd_sc_hd__a21o_1
Xhold556 la_data_in[30] vssd2 vssd2 vccd2 vccd2 hold49/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 input45/X vssd2 vssd2 vccd2 vccd2 hold82/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold567 hold66/X vssd2 vssd2 vccd2 vccd2 _7860_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_474 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_40_485 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold589 hold87/X vssd2 vssd2 vccd2 vccd2 input44/A sky130_fd_sc_hd__dlygate4sd3_1
X_6225_ _6221_/X _6223_/X _6152_/B vssd2 vssd2 vccd2 vccd2 _7140_/A sky130_fd_sc_hd__o21ai_4
XTAP_861 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _6154_/Y _6155_/X _6100_/D _6587_/B _5938_/C vssd2 vssd2 vccd2 vccd2 _6156_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_894 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _5178_/B _5107_/B vssd2 vssd2 vccd2 vccd2 _5110_/A sky130_fd_sc_hd__nor2_2
X_6087_ _6707_/A _6581_/A vssd2 vssd2 vccd2 vccd2 _6091_/A sky130_fd_sc_hd__nor2_1
X_5038_ _5052_/A vssd2 vssd2 vccd2 vccd2 _5038_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_79_165 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_79_187 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6989_ _6989_/A _7255_/B vssd2 vssd2 vccd2 vccd2 _6991_/B sky130_fd_sc_hd__nor2_1
XANTENNA__6935__A2 _6040_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_82_319 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_63_544 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_63_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_63_599 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_105_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_50_249 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4174__A2 _4044_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_98_441 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_85_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_39_530 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_160 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_54_511 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_39_585 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_193 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_182 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_171 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6033__B _6855_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_54_555 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_54_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_109_495 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_41_249 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7145__A _7145_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_111_137 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4340_ _4277_/A _4276_/A _4276_/B vssd2 vssd2 vccd2 vccd2 _4347_/A sky130_fd_sc_hd__a21boi_4
X_4271_ _4266_/X _4270_/X _3996_/B vssd2 vssd2 vccd2 vccd2 _4271_/Y sky130_fd_sc_hd__o21ai_1
X_6010_ _6064_/B _6010_/B vssd2 vssd2 vccd2 vccd2 _6068_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_441 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6912_ _7033_/A _7033_/B _7033_/C _7034_/A vssd2 vssd2 vccd2 vccd2 _6970_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_89_474 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_49_305 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6843_ _6909_/B _6843_/B vssd2 vssd2 vccd2 vccd2 _7824_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_76_135 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__3848__A _4267_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_91_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4928__A1 _4863_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6774_ _6776_/A _6776_/B _6776_/C vssd2 vssd2 vccd2 vccd2 _6901_/A sky130_fd_sc_hd__a21oi_2
X_3986_ _3986_/A _3986_/B vssd2 vssd2 vccd2 vccd2 _3986_/X sky130_fd_sc_hd__and2_1
XFILLER_0_91_149 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_84_190 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_57_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5725_ _6152_/B _5944_/B _5937_/B _5769_/B vssd2 vssd2 vccd2 vccd2 _5845_/C sky130_fd_sc_hd__or4_1
XFILLER_0_94_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_72_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5656_ _5653_/X _5655_/X _6396_/B vssd2 vssd2 vccd2 vccd2 _5674_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_72_396 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4607_ _4535_/A _4535_/B _4533_/X vssd2 vssd2 vccd2 vccd2 _4609_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_60_569 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5587_ _5583_/A _5583_/B _5586_/Y vssd2 vssd2 vccd2 vccd2 _5587_/X sky130_fd_sc_hd__a21o_1
Xhold320 _7485_/X vssd2 vssd2 vccd2 vccd2 _7725_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_290 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7326_ _7326_/A _7326_/B _7326_/C _7326_/D vssd2 vssd2 vccd2 vccd2 _7335_/B sky130_fd_sc_hd__nand4_2
X_4538_ _4538_/A _4538_/B vssd2 vssd2 vccd2 vccd2 _4539_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__4398__B _4966_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold353 _7754_/Q vssd2 vssd2 vccd2 vccd2 hold353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 _7477_/X vssd2 vssd2 vccd2 vccd2 _7717_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 _7745_/Q vssd2 vssd2 vccd2 vccd2 hold331/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_496 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7257_ _7181_/A _6670_/Y _7256_/Y vssd2 vssd2 vccd2 vccd2 _7259_/C sky130_fd_sc_hd__o21a_1
X_4469_ _4469_/A _4469_/B vssd2 vssd2 vccd2 vccd2 _4470_/B sky130_fd_sc_hd__xor2_4
Xhold364 _7691_/Q vssd2 vssd2 vccd2 vccd2 hold364/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_94 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold375 _7650_/Q vssd2 vssd2 vccd2 vccd2 hold375/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 _7684_/Q vssd2 vssd2 vccd2 vccd2 hold386/X sky130_fd_sc_hd__dlygate4sd3_1
X_6208_ _6208_/A _6208_/B vssd2 vssd2 vccd2 vccd2 _6210_/B sky130_fd_sc_hd__xnor2_2
Xhold397 hold693/X vssd2 vssd2 vccd2 vccd2 _7770_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7188_ _7188_/A _7188_/B vssd2 vssd2 vccd2 vccd2 _7189_/B sky130_fd_sc_hd__or2_1
XFILLER_0_99_205 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6139_ _6139_/A _6139_/B vssd2 vssd2 vccd2 vccd2 _6140_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__5408__A2 _5550_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_680 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_249 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4564__D _4782_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_68_614 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_67_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_95_444 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4861__B _5168_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5041__B1 _5528_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_75_190 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_36_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__5973__A _6138_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4589__A _4810_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_31_260 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_48_17 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_101_181 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6028__B _6783_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_80_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_58_146 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_86_488 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_13_31 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_13_42 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_3840_ _3813_/A _3813_/B _4458_/D _4144_/C _4326_/C vssd2 vssd2 vccd2 vccd2 _4141_/C
+ sky130_fd_sc_hd__a2111o_2
XFILLER_0_104_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6780__B1 _7222_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_6_405 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_109_281 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_42_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5510_ _5510_/A _5510_/B vssd2 vssd2 vccd2 vccd2 _5512_/B sky130_fd_sc_hd__xnor2_1
X_6490_ _6491_/B _6491_/A vssd2 vssd2 vccd2 vccd2 _6490_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_89_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_112_413 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5441_ _5392_/A _5392_/B _5393_/X vssd2 vssd2 vccd2 vccd2 _5443_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_42_569 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_112_457 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5372_ _5330_/A _5330_/B _5329_/B vssd2 vssd2 vccd2 vccd2 _5377_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__7088__B2 _6571_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7111_ _7111_/A _7111_/B vssd2 vssd2 vccd2 vccd2 _7117_/A sky130_fd_sc_hd__xor2_1
X_4323_ _4323_/A _4323_/B _4323_/C vssd2 vssd2 vccd2 vccd2 _4324_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_1_176 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7042_ _7042_/A _7042_/B vssd2 vssd2 vccd2 vccd2 _7064_/A sky130_fd_sc_hd__xor2_1
XANTENNA__7603__A _7627_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4254_ _4252_/X _4253_/Y _4707_/A vssd2 vssd2 vccd2 vccd2 _4254_/Y sky130_fd_sc_hd__a21oi_1
X_4185_ _4186_/A _4186_/B vssd2 vssd2 vccd2 vccd2 _4243_/A sky130_fd_sc_hd__or2_1
XANTENNA__4962__A _4962_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_89_293 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_77_422 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1109 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4074__B2 _4162_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4074__A1 _7768_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_fanout265_A _7848_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7875_ _7878_/CLK _7875_/D _7634_/Y vssd2 vssd2 vccd2 vccd2 _7875_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_499 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6826_ _6826_/A _6826_/B vssd2 vssd2 vccd2 vccd2 _6829_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_617 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_64_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6757_ _6757_/A _6757_/B vssd2 vssd2 vccd2 vccd2 _6758_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_149 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_64_127 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_18_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5708_ _5694_/A _5694_/B _5735_/B vssd2 vssd2 vccd2 vccd2 _5711_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_9_298 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3969_ _3967_/X _3968_/X _3943_/X vssd2 vssd2 vccd2 vccd2 _3969_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_33_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6688_ _6688_/A _6688_/B vssd2 vssd2 vccd2 vccd2 _6689_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_72_171 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_33_525 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6401__B _7253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5639_ _7856_/Q _7855_/Q _7857_/Q _5645_/B vssd2 vssd2 vccd2 vccd2 _5640_/B sky130_fd_sc_hd__o31a_2
XFILLER_0_79_90 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4202__A _7768_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_103_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7309_ _7309_/A _7309_/B vssd2 vssd2 vccd2 vccd2 _7326_/D sky130_fd_sc_hd__xnor2_2
Xhold150 hold360/X vssd2 vssd2 vccd2 vccd2 _7790_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 _7388_/X vssd2 vssd2 vccd2 vccd2 _7389_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7513__A _7641_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold183 _7365_/X vssd2 vssd2 vccd2 vccd2 _7366_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 input87/X vssd2 vssd2 vccd2 vccd2 hold194/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 input94/X vssd2 vssd2 vccd2 vccd2 hold172/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_6 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1632 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_455 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_68_499 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_68_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_55_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_83_469 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_71_609 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7394__S _7418_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_36_352 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_525 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_75_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_99_591 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4782__A _5210_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_400 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5990_ _7847_/Q _6357_/B _5989_/X _5944_/C vssd2 vssd2 vccd2 vccd2 _5990_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_91_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4941_ _4941_/A _4941_/B vssd2 vssd2 vccd2 vccd2 _4943_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_444 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4872_ _4872_/A _4872_/B vssd2 vssd2 vccd2 vccd2 _4873_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_116 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7660_ _7806_/CLK _7660_/D vssd2 vssd2 vccd2 vccd2 _7660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_52 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6611_ _6694_/A _6611_/B vssd2 vssd2 vccd2 vccd2 _6613_/B sky130_fd_sc_hd__and2_1
XFILLER_0_46_127 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3823_ _3822_/A _3822_/B _3822_/C _3821_/X _3888_/B vssd2 vssd2 vccd2 vccd2 _3825_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_0_24_96 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7591_ _7597_/A vssd2 vssd2 vccd2 vccd2 _7591_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4006__B _4006_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6542_ _6542_/A _6542_/B vssd2 vssd2 vccd2 vccd2 _6608_/A sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_9_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7758_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_525 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6473_ _6474_/A _6474_/B vssd2 vssd2 vccd2 vccd2 _7222_/C sky130_fd_sc_hd__and2_4
XFILLER_0_42_355 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_112_221 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5424_ _5424_/A _5424_/B vssd2 vssd2 vccd2 vccd2 _5427_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_112_265 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_100_416 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_42_399 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_2_474 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7333__A _7333_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5355_ _5254_/A _5254_/B _5308_/A _5354_/X vssd2 vssd2 vccd2 vccd2 _5356_/B sky130_fd_sc_hd__a31o_2
XFILLER_0_57_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5286_ _5287_/A _5287_/B vssd2 vssd2 vccd2 vccd2 _5341_/B sky130_fd_sc_hd__and2b_1
X_4306_ _5548_/A _4308_/B vssd2 vssd2 vccd2 vccd2 _4307_/B sky130_fd_sc_hd__nor2_1
X_7025_ _7025_/A _7025_/B _7025_/C _7025_/D vssd2 vssd2 vccd2 vccd2 _7025_/X sky130_fd_sc_hd__or4_2
X_4237_ _4237_/A _4237_/B vssd2 vssd2 vccd2 vccd2 _4239_/A sky130_fd_sc_hd__xor2_1
X_4168_ _7765_/Q _4814_/B _4707_/A vssd2 vssd2 vccd2 vccd2 _4168_/X sky130_fd_sc_hd__and3_1
XFILLER_0_97_528 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4099_ _7765_/Q _4454_/B vssd2 vssd2 vccd2 vccd2 _4099_/X sky130_fd_sc_hd__and2_1
X_7858_ _7886_/CLK _7858_/D _7617_/Y vssd2 vssd2 vccd2 vccd2 _7858_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_92_233 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6809_ _6808_/B _6808_/C _6808_/A vssd2 vssd2 vccd2 vccd2 _6820_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_277 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7789_ _7806_/CLK _7789_/D _7548_/Y vssd2 vssd2 vccd2 vccd2 _7789_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_80_439 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_333 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_60_152 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__5028__A _5029_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_21_517 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5786__A1 _7846_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1440 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_414 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5210__B _5210_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_29_617 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1484 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_211 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_68_296 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_56_425 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1495 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6735__B1 _7222_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_43_108 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_71_428 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_9_18 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4210__A1 _4328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_64_491 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_344 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_355 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4210__B2 _7767_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_51_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_10_32 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_12_506 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_377 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6976__B _7291_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4777__A _4863_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4496__B _4896_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5140_ _5011_/A _5431_/B _5243_/A _5139_/X vssd2 vssd2 vccd2 vccd2 _5187_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_20_583 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5071_ _5072_/A _5072_/B _5072_/C vssd2 vssd2 vccd2 vccd2 _5192_/A sky130_fd_sc_hd__o21a_2
X_4022_ _4315_/B _4022_/B _4427_/A vssd2 vssd2 vccd2 vccd2 _4160_/B sky130_fd_sc_hd__and3_2
X_5973_ _6138_/A _6812_/A vssd2 vssd2 vccd2 vccd2 _5974_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5777__A1 _6158_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4924_ _4924_/A _4924_/B vssd2 vssd2 vccd2 vccd2 _4925_/B sky130_fd_sc_hd__nor2_2
XANTENNA__4662__D _5315_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_274 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7712_ _7771_/CLK _7712_/D vssd2 vssd2 vccd2 vccd2 _7712_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5777__B2 _6157_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_74_222 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_47_425 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4855_ _4990_/A _4855_/B vssd2 vssd2 vccd2 vccd2 _4855_/Y sky130_fd_sc_hd__nand2b_1
X_7643_ _7645_/A vssd2 vssd2 vccd2 vccd2 _7643_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_661 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7328__A _7334_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7574_ _7613_/A vssd2 vssd2 vccd2 vccd2 _7574_/Y sky130_fd_sc_hd__inv_2
X_4786_ _4714_/A _4714_/B _4712_/B vssd2 vssd2 vccd2 vccd2 _4787_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_62_417 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3806_ _7793_/Q _7792_/Q _7791_/Q _7794_/Q vssd2 vssd2 vccd2 vccd2 _3822_/A sky130_fd_sc_hd__or4_4
XFILLER_0_34_108 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6525_ _6446_/A _6446_/B _6444_/X vssd2 vssd2 vccd2 vccd2 _6527_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_113_541 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_15_355 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_30_303 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_42_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6456_ _6457_/A _6457_/B vssd2 vssd2 vccd2 vccd2 _6456_/Y sky130_fd_sc_hd__nor2_1
X_6387_ _6387_/A _6387_/B _6387_/C vssd2 vssd2 vccd2 vccd2 _6387_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_11_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5407_ _5407_/A _5407_/B vssd2 vssd2 vccd2 vccd2 _5407_/Y sky130_fd_sc_hd__xnor2_1
X_5338_ _5339_/B _5339_/A vssd2 vssd2 vccd2 vccd2 _5338_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_2_293 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7008_ _6939_/A _7255_/B _6940_/A _6937_/X vssd2 vssd2 vccd2 vccd2 _7008_/X sky130_fd_sc_hd__o31a_1
X_5269_ _5270_/A _5270_/B vssd2 vssd2 vccd2 vccd2 _5379_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__5014__C _5414_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_78_550 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5030__B _5030_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_65_233 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_38_447 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_53_406 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_108_357 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_65_299 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_65_277 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6193__A1 _7849_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_46_491 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6193__B2 _7850_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4743__A2 _4809_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7142__B1 _7313_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3951__B1 _4050_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_33_185 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XTAP_509 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5205__B _5404_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout290 _7597_/A vssd2 vssd2 vccd2 vccd2 _7590_/A sky130_fd_sc_hd__buf_8
XANTENNA__6317__A _7034_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_69_572 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1292 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_233 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_84_586 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4640_ _4640_/A _4640_/B vssd2 vssd2 vccd2 vccd2 _4641_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_417 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_21_31 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_114_305 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_112_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_71_236 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_37_491 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_114_349 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6310_ _6387_/B _6310_/B vssd2 vssd2 vccd2 vccd2 _6313_/A sky130_fd_sc_hd__xnor2_1
X_4571_ _4572_/A _4572_/B vssd2 vssd2 vccd2 vccd2 _4571_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__6987__A _7045_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5891__A _6424_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_24_163 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7290_ _7319_/A _7290_/B vssd2 vssd2 vccd2 vccd2 _7297_/A sky130_fd_sc_hd__and2_1
XFILLER_0_40_645 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_110_533 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6241_ _6241_/A _6241_/B vssd2 vssd2 vccd2 vccd2 _6242_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6172_ _6172_/A _6172_/B vssd2 vssd2 vccd2 vccd2 _6173_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_110_577 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5123_ _5123_/A _5123_/B vssd2 vssd2 vccd2 vccd2 _5126_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__7611__A _7613_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5054_ _5055_/B _5055_/A vssd2 vssd2 vccd2 vccd2 _5054_/X sky130_fd_sc_hd__and2b_1
XANTENNA__4954__B _5030_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4005_ _7765_/Q _4458_/D _4268_/D vssd2 vssd2 vccd2 vccd2 _4005_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_79_358 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5956_ _5956_/A _5956_/B _5956_/C vssd2 vssd2 vccd2 vccd2 _5958_/B sky130_fd_sc_hd__or3_1
XFILLER_0_75_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4907_ _4907_/A _4907_/B vssd2 vssd2 vccd2 vccd2 _4908_/B sky130_fd_sc_hd__xor2_4
X_5887_ _5885_/X _5886_/X _6424_/A vssd2 vssd2 vccd2 vccd2 _5890_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_90_501 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4838_ _4839_/A _4839_/B vssd2 vssd2 vccd2 vccd2 _4923_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_62_214 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7626_ _7627_/A vssd2 vssd2 vccd2 vccd2 _7626_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_105_305 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_105_349 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4769_ _4769_/A _4769_/B vssd2 vssd2 vccd2 vccd2 _7740_/D sky130_fd_sc_hd__xnor2_2
X_7557_ _7557_/A vssd2 vssd2 vccd2 vccd2 _7557_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5009__C _5142_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6508_ _6668_/A _7099_/B vssd2 vssd2 vccd2 vccd2 _6516_/A sky130_fd_sc_hd__nand2_1
X_7488_ _7524_/A vssd2 vssd2 vccd2 vccd2 _7488_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3933__B1 _4050_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_101_511 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__6478__A2 _6404_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6439_ _6668_/A _7197_/A _6365_/B _6363_/X vssd2 vssd2 vccd2 vccd2 _6441_/B sky130_fd_sc_hd__a31o_1
XANTENNA__5951__D _6855_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_113_393 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_101_599 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xhold32 hold32/A vssd2 vssd2 vccd2 vccd2 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd2 vssd2 vccd2 vccd2 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd2 vssd2 vccd2 vccd2 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7521__A _7557_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold43 hold43/A vssd2 vssd2 vccd2 vccd2 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5989__A1 _6158_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5989__B2 _6283_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold65 hold65/A vssd2 vssd2 vccd2 vccd2 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd2 vssd2 vccd2 vccd2 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd2 vssd2 vccd2 vccd2 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd2 vssd2 vccd2 vccd2 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd2 vssd2 vccd2 vccd2 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4661__B2 _4807_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_85_328 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_66_520 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4880__A _5029_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_38_244 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_108_121 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_66_597 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_108_165 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7115__B1 _7047_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_7 hold84/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_22_623 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_22_645 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_104_371 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_21_122 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_306 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4120__A _4656_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5141__A2 _5142_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_339 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6973__C _7253_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_83_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_wb_clk_i clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7793_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_107_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_89_645 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_88_166 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_49_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6790_ _6790_/A _6790_/B vssd2 vssd2 vccd2 vccd2 _6793_/A sky130_fd_sc_hd__nand2_1
X_5810_ _6016_/B _6071_/B vssd2 vssd2 vccd2 vccd2 _5810_/X sky130_fd_sc_hd__and2_1
X_5741_ _5769_/B _5992_/B vssd2 vssd2 vccd2 vccd2 _5742_/D sky130_fd_sc_hd__nor2_1
XANTENNA__5601__B1 _5645_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_84_361 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_84_350 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4940__D _5315_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_8_149 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_32_52 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7411_ _7452_/A _7411_/B vssd2 vssd2 vccd2 vccd2 _7411_/X sky130_fd_sc_hd__and2_1
X_5672_ _5650_/X _5671_/X _5670_/X vssd2 vssd2 vccd2 vccd2 _5672_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_32_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_114_113 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_72_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_72_578 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4623_ _4614_/A _4614_/B _4612_/Y vssd2 vssd2 vccd2 vccd2 _4683_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_25_461 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_32_409 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7606__A _7627_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3915__B1 _4050_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7342_ _7342_/A _7342_/B _7342_/C _7342_/D vssd2 vssd2 vccd2 vccd2 _7345_/B sky130_fd_sc_hd__or4_1
X_4554_ _5455_/A _4556_/B vssd2 vssd2 vccd2 vccd2 _4555_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_13_634 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold502 input20/X vssd2 vssd2 vccd2 vccd2 hold48/A sky130_fd_sc_hd__dlygate4sd3_1
X_7273_ _7273_/A _7273_/B vssd2 vssd2 vccd2 vccd2 _7274_/B sky130_fd_sc_hd__and2_1
Xhold524 la_data_in[23] vssd2 vssd2 vccd2 vccd2 hold59/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold535 hold58/X vssd2 vssd2 vccd2 vccd2 _7864_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 hold45/X vssd2 vssd2 vccd2 vccd2 input19/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 input40/X vssd2 vssd2 vccd2 vccd2 hold70/A sky130_fd_sc_hd__dlygate4sd3_1
X_4485_ _4475_/A _4475_/B _4473_/Y vssd2 vssd2 vccd2 vccd2 _4545_/A sky130_fd_sc_hd__a21boi_2
Xhold557 hold49/X vssd2 vssd2 vccd2 vccd2 input24/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_188 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold579 hold82/X vssd2 vssd2 vccd2 vccd2 _7877_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 la_data_in[16] vssd2 vssd2 vccd2 vccd2 hold85/A sky130_fd_sc_hd__dlygate4sd3_1
X_6224_ _6221_/X _6223_/X _6152_/B vssd2 vssd2 vccd2 vccd2 _7197_/A sky130_fd_sc_hd__o21a_4
XFILLER_0_110_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4965__A _5220_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_862 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _6152_/B _6155_/B _6253_/A vssd2 vssd2 vccd2 vccd2 _6155_/X sky130_fd_sc_hd__and3b_1
X_6086_ _6086_/A _6086_/B vssd2 vssd2 vccd2 vccd2 _6115_/A sky130_fd_sc_hd__xnor2_1
XTAP_895 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4891__B2 _4962_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_873 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _5164_/A _5105_/B _5105_/C vssd2 vssd2 vccd2 vccd2 _5107_/B sky130_fd_sc_hd__o21a_1
X_5037_ _5091_/B _5037_/B vssd2 vssd2 vccd2 vccd2 _5052_/A sky130_fd_sc_hd__or2_2
XFILLER_0_73_81 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__5199__A2 _5528_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_82_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6988_ _6988_/A _6988_/B vssd2 vssd2 vccd2 vccd2 _6991_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_542 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6404__B _6634_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_75_350 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5939_ _7844_/Q _6510_/B vssd2 vssd2 vccd2 vccd2 _5939_/X sky130_fd_sc_hd__and2_1
XFILLER_0_63_556 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_35_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_247 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_105_113 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7609_ _7613_/A vssd2 vssd2 vccd2 vccd2 _7609_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7516__A _7564_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_16_472 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_31_486 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_101_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_9_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xinput100 wbs_we_i vssd2 vssd2 vccd2 vccd2 _7350_/C sky130_fd_sc_hd__buf_1
XFILLER_0_98_453 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_86_648 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_39_520 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_542 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_39_553 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_85_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XPHY_161 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_150 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_66_361 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_109_452 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_194 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_183 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_172 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_26_247 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6330__A _6402_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_81_397 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_81_386 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_78_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__3954__A _4050_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7426__A _7436_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_111_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__7145__B _7222_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4769__B _4769_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_34_291 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_111_149 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4270_ _4454_/A _4075_/B _4267_/X _4268_/X _4269_/X vssd2 vssd2 vccd2 vccd2 _4270_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__5822__B1 _7336_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6911_ _7033_/B _6911_/B vssd2 vssd2 vccd2 vccd2 _7825_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_77_615 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_77_604 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6842_ _6909_/A _7033_/A _7034_/A vssd2 vssd2 vccd2 vccd2 _6843_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_43_62 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4928__A2 _5550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6773_ _6707_/A _6549_/Y _6704_/X _6706_/B vssd2 vssd2 vccd2 vccd2 _6776_/C sky130_fd_sc_hd__o31a_1
XFILLER_0_64_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_9_447 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3985_ _4214_/C _4018_/A _4164_/C _5030_/A vssd2 vssd2 vccd2 vccd2 _3986_/B sky130_fd_sc_hd__nor4_1
XANTENNA__7327__B1 _6069_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5724_ _6152_/B _5944_/B _5937_/B _5769_/B vssd2 vssd2 vccd2 vccd2 _5898_/C sky130_fd_sc_hd__nor4_1
XFILLER_0_17_236 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_45_556 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_17_269 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5655_ _6253_/B _5655_/B _5655_/C vssd2 vssd2 vccd2 vccd2 _5655_/X sky130_fd_sc_hd__and3_1
XFILLER_0_32_206 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7336__A _7336_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4606_ _4606_/A _4606_/B vssd2 vssd2 vccd2 vccd2 _4609_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_526 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5889__B1 _6424_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7325_ _7334_/C vssd2 vssd2 vccd2 vccd2 _7325_/Y sky130_fd_sc_hd__inv_2
Xhold310 hold310/A vssd2 vssd2 vccd2 vccd2 la_data_out[24] sky130_fd_sc_hd__buf_12
X_5586_ _7870_/Q _5586_/B vssd2 vssd2 vccd2 vccd2 _5586_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_13_431 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4537_ _4538_/A _4538_/B vssd2 vssd2 vccd2 vccd2 _4537_/Y sky130_fd_sc_hd__nand2b_1
Xhold321 _7756_/Q vssd2 vssd2 vccd2 vccd2 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 _7750_/Q vssd2 vssd2 vccd2 vccd2 hold343/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 _7473_/X vssd2 vssd2 vccd2 vccd2 _7713_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_464 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4468_ _4468_/A _4468_/B vssd2 vssd2 vccd2 vccd2 _4469_/B sky130_fd_sc_hd__xnor2_2
X_7256_ _7256_/A _7256_/B vssd2 vssd2 vccd2 vccd2 _7256_/Y sky130_fd_sc_hd__xnor2_1
Xhold387 _7657_/Q vssd2 vssd2 vccd2 vccd2 hold387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 hold686/X vssd2 vssd2 vccd2 vccd2 _7797_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 hold682/X vssd2 vssd2 vccd2 vccd2 _7783_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 _7482_/X vssd2 vssd2 vccd2 vccd2 _7722_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6207_ _6636_/A _7037_/A _6208_/B vssd2 vssd2 vccd2 vccd2 _6207_/X sky130_fd_sc_hd__or3_1
X_7187_ _7188_/A _7188_/B vssd2 vssd2 vccd2 vccd2 _7232_/B sky130_fd_sc_hd__nand2_1
Xhold398 hold695/X vssd2 vssd2 vccd2 vccd2 _7774_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4695__A _5548_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6138_ _6138_/A _6973_/A vssd2 vssd2 vccd2 vccd2 _6139_/B sky130_fd_sc_hd__nor2_1
X_4399_ wire212/X _4881_/A2 _5099_/A vssd2 vssd2 vccd2 vccd2 _4401_/B sky130_fd_sc_hd__a21oi_2
XTAP_670 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6066__B1 _7336_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_681 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _6069_/A _6189_/A vssd2 vssd2 vccd2 vccd2 _6127_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_95_412 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_95_401 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_68_648 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4861__C _5142_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_67_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5041__A1 _5145_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5041__B2 _5042_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_36_501 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5973__B _6812_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_106_455 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6150__A _6150_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_63_375 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6788__C _7181_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4589__B _5406_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_31_272 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_101_193 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5804__B1 _7843_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_80_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_73_117 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_46_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6780__A1 _5994_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_54_331 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_6_417 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_13_65 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6780__B2 _5948_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_13_76 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_109_293 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_54_386 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_42_537 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_42_526 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5440_ _5486_/B _5440_/B vssd2 vssd2 vccd2 vccd2 _5443_/A sky130_fd_sc_hd__and2_1
XFILLER_0_89_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_1_100 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5371_ _5430_/A _5371_/B vssd2 vssd2 vccd2 vccd2 _5382_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_112_469 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__7088__A2 _7313_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7110_ _7111_/A _7111_/B vssd2 vssd2 vccd2 vccd2 _7166_/A sky130_fd_sc_hd__nor2_1
X_4322_ _4323_/A _4323_/B _4323_/C vssd2 vssd2 vccd2 vccd2 _4413_/A sky130_fd_sc_hd__o21a_2
X_7041_ _7040_/A _7040_/B _7042_/A vssd2 vssd2 vccd2 vccd2 _7106_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_59_7 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4253_ _7768_/Q _4253_/B vssd2 vssd2 vccd2 vccd2 _4253_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5404__A _5404_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4184_ _4136_/A _4136_/B _4135_/A vssd2 vssd2 vccd2 vccd2 _4186_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_38_95 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_96_209 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_89_261 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA_fanout258_A _7853_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7874_ _7878_/CLK _7874_/D _7633_/Y vssd2 vssd2 vccd2 vccd2 _7874_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_478 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6825_ _6825_/A _6825_/B vssd2 vssd2 vccd2 vccd2 _6826_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_117 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_49_158 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_9_222 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6756_ _6757_/A _6757_/B vssd2 vssd2 vccd2 vccd2 _6756_/X sky130_fd_sc_hd__or2_1
XFILLER_0_64_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3968_ _4022_/B _4162_/B _7766_/Q vssd2 vssd2 vccd2 vccd2 _3968_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_45_364 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_18_556 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5707_ _6283_/B _6094_/B _6510_/B _6670_/B vssd2 vssd2 vccd2 vccd2 _6102_/B sky130_fd_sc_hd__nor4_4
X_6687_ _6688_/A _6688_/B vssd2 vssd2 vccd2 vccd2 _6687_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_60_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_3899_ _7791_/Q _7768_/Q _4006_/C _3899_/D vssd2 vssd2 vccd2 vccd2 _3899_/X sky130_fd_sc_hd__and4_1
XFILLER_0_72_194 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5638_ _6158_/A _5638_/B _5638_/C vssd2 vssd2 vccd2 vccd2 _5638_/X sky130_fd_sc_hd__and3_1
XFILLER_0_33_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5569_ _5556_/A _5556_/B _5568_/Y vssd2 vssd2 vccd2 vccd2 _5570_/C sky130_fd_sc_hd__o21ai_1
X_7308_ _7308_/A _7308_/B vssd2 vssd2 vccd2 vccd2 _7309_/B sky130_fd_sc_hd__nand2_1
Xhold151 _7418_/X vssd2 vssd2 vccd2 vccd2 _7419_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 hold364/X vssd2 vssd2 vccd2 vccd2 _7803_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 _7435_/X vssd2 vssd2 vccd2 vccd2 _7436_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_592 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold173 _7398_/X vssd2 vssd2 vccd2 vccd2 _7399_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _7414_/X vssd2 vssd2 vccd2 vccd2 _7415_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 hold380/X vssd2 vssd2 vccd2 vccd2 _7764_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7239_ _7239_/A _7239_/B _7239_/C vssd2 vssd2 vccd2 vccd2 _7240_/B sky130_fd_sc_hd__or3_1
XTAP_1600 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6145__A _6634_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_68_434 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4591__C _5042_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_83_404 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_68_489 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_49_670 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_28_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_83_437 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5984__A _6550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_117 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_50_19 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_36_397 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_63_194 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_51_345 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_59_17 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_51_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_75_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_91_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5253__A1 _4996_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4782__B _4782_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_231 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4940_ _5210_/A _5210_/B _5222_/A _5315_/B vssd2 vssd2 vccd2 vccd2 _4941_/B sky130_fd_sc_hd__or4_1
XFILLER_0_86_253 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4871_ _4872_/A _4872_/B vssd2 vssd2 vccd2 vccd2 _4873_/A sky130_fd_sc_hd__or2_1
XFILLER_0_59_467 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__3829__D _4006_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7590_ _7590_/A vssd2 vssd2 vccd2 vccd2 _7590_/Y sky130_fd_sc_hd__inv_2
X_6610_ _6610_/A _6610_/B _6610_/C vssd2 vssd2 vccd2 vccd2 _6611_/B sky130_fd_sc_hd__nand3_1
X_3822_ _3822_/A _3822_/B _3822_/C _3822_/D vssd2 vssd2 vccd2 vccd2 _3822_/X sky130_fd_sc_hd__or4_1
XFILLER_0_27_320 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6541_ _6542_/A _6542_/B vssd2 vssd2 vccd2 vccd2 _6693_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_74_459 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_109 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_54_194 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6472_ _6398_/A _7313_/A _6194_/B _6670_/A vssd2 vssd2 vccd2 vccd2 _6474_/B sky130_fd_sc_hd__a22o_2
XFILLER_0_15_548 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_40_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_112_233 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_30_529 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5423_ _5424_/A _5424_/B vssd2 vssd2 vccd2 vccd2 _5472_/B sky130_fd_sc_hd__nor2_1
X_5354_ _5247_/A _5303_/Y _5304_/Y vssd2 vssd2 vccd2 vccd2 _5354_/X sky130_fd_sc_hd__o21a_1
XANTENNA__7614__A _7641_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_112_277 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_49_61 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4305_ _4305_/A _4305_/B vssd2 vssd2 vccd2 vccd2 _4308_/B sky130_fd_sc_hd__and2_1
X_5285_ _5328_/A _5550_/A vssd2 vssd2 vccd2 vccd2 _5287_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5134__A _5455_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7024_ _7024_/A _7024_/B vssd2 vssd2 vccd2 vccd2 _7211_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__7481__A2 _7483_/A2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4236_ _4237_/A _4237_/B vssd2 vssd2 vccd2 vccd2 _4236_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4167_ _4161_/Y _4166_/X _4125_/C vssd2 vssd2 vccd2 vccd2 _4171_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_97_518 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4098_ _4898_/A _4807_/A vssd2 vssd2 vccd2 vccd2 _4118_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_77_231 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7857_ _7886_/CLK _7857_/D _7616_/Y vssd2 vssd2 vccd2 vccd2 _7857_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_65_437 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6808_ _6808_/A _6808_/B _6808_/C vssd2 vssd2 vccd2 vccd2 _6820_/A sky130_fd_sc_hd__and3_1
XFILLER_0_92_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7788_ _7806_/CLK _7788_/D _7547_/Y vssd2 vssd2 vccd2 vccd2 _7788_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_92_289 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_73_481 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6739_ _6739_/A _6739_/B vssd2 vssd2 vccd2 vccd2 _6742_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_60_131 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_33_345 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_61_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_60_164 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_33_367 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7472__A2 _7483_/A2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5979__A _6670_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1441 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_573 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_96_551 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_68_253 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5210__C _5528_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1474 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_448 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1496 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6735__B2 _6664_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6735__A1 _6424_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_107_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_3_206 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_101_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7160__A1 _7045_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7434__A _7436_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4777__B _5011_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4496__C _4711_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5070_ _5008_/X _5012_/B _5010_/B vssd2 vssd2 vccd2 vccd2 _5072_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__7463__A2 _7454_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6671__B1 _6669_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4021_ _4328_/A _4214_/C _4125_/C _4021_/D vssd2 vssd2 vccd2 vccd2 _4021_/X sky130_fd_sc_hd__and4_1
X_5972_ _5778_/X _5786_/Y _6812_/B _5736_/X vssd2 vssd2 vccd2 vccd2 _5974_/A sky130_fd_sc_hd__a211o_1
XFILLER_0_59_231 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5777__A2 _5992_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4923_ _4923_/A _4923_/B _4923_/C vssd2 vssd2 vccd2 vccd2 _4924_/B sky130_fd_sc_hd__and3_1
X_7711_ _7771_/CLK _7711_/D vssd2 vssd2 vccd2 vccd2 _7711_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__7609__A _7613_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_47_437 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_4854_ _4854_/A _4854_/B _4854_/C vssd2 vssd2 vccd2 vccd2 _4855_/B sky130_fd_sc_hd__or3_1
X_7642_ _7645_/A vssd2 vssd2 vccd2 vccd2 _7642_/Y sky130_fd_sc_hd__inv_2
X_7573_ _7613_/A vssd2 vssd2 vccd2 vccd2 _7573_/Y sky130_fd_sc_hd__inv_2
X_4785_ _4785_/A _4785_/B vssd2 vssd2 vccd2 vccd2 _4787_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_62_429 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3805_ _7524_/A vssd2 vssd2 vccd2 vccd2 _7450_/A sky130_fd_sc_hd__inv_2
X_6524_ _6524_/A _6524_/B vssd2 vssd2 vccd2 vccd2 _6527_/A sky130_fd_sc_hd__xor2_2
XANTENNA__4033__A _7768_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_43_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_113_553 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6455_ _6455_/A _6455_/B vssd2 vssd2 vccd2 vccd2 _6457_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_175 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_42_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6386_ _6387_/A _6387_/B _6387_/C vssd2 vssd2 vccd2 vccd2 _6389_/A sky130_fd_sc_hd__and3_1
X_5406_ _5406_/A _5550_/A vssd2 vssd2 vccd2 vccd2 _5407_/B sky130_fd_sc_hd__nor2_1
X_5337_ _5293_/A _5293_/B _5274_/Y vssd2 vssd2 vccd2 vccd2 _5339_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_76_70 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5268_ _5225_/A _5225_/B _5223_/Y vssd2 vssd2 vccd2 vccd2 _5270_/B sky130_fd_sc_hd__o21ai_2
X_7007_ _7007_/A _7007_/B _7007_/C vssd2 vssd2 vccd2 vccd2 _7012_/B sky130_fd_sc_hd__and3_1
X_4219_ _4598_/A _4219_/B _4662_/B vssd2 vssd2 vccd2 vccd2 _4220_/B sky130_fd_sc_hd__or3_1
XANTENNA__5014__D _5081_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5199_ _4172_/Y _5528_/A _5029_/X _5160_/B _5163_/A vssd2 vssd2 vccd2 vccd2 _5201_/C
+ sky130_fd_sc_hd__o41a_1
XANTENNA__5762__A_N _5736_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4208__A _4810_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_78_562 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_93_510 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_78_595 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7519__A _7557_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6423__A _6425_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_38_459 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_53_418 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_46_481 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_61_495 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_484 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__7142__A1 _7143_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7142__B2 _7143_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_21_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_104_575 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5205__C _5414_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout291 _7629_/A vssd2 vssd2 vccd2 vccd2 _7597_/A sky130_fd_sc_hd__buf_4
Xfanout280 _7450_/A vssd2 vssd2 vccd2 vccd2 _7452_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_551 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_84_521 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_69_584 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__4967__B1 _5528_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_8_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XTAP_1293 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4570_ _4570_/A _4570_/B vssd2 vssd2 vccd2 vccd2 _4572_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_108_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_107_391 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6987__B _7253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_12_304 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6240_ _6241_/B _6241_/A vssd2 vssd2 vccd2 vccd2 _6240_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_97_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_12_359 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_110_545 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6171_ _6172_/A _6172_/B vssd2 vssd2 vccd2 vccd2 _6171_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_110_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5122_ _5122_/A _5122_/B vssd2 vssd2 vccd2 vccd2 _5123_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__6508__A _6668_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5053_ _4978_/A _4978_/B _4976_/Y vssd2 vssd2 vccd2 vccd2 _5055_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_46_62 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4004_ _4454_/A _4004_/B vssd2 vssd2 vccd2 vccd2 _4004_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_94_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5955_ _5956_/A _5956_/B _5956_/C vssd2 vssd2 vccd2 vccd2 _5955_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_47_212 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4906_ _4907_/A _4907_/B vssd2 vssd2 vccd2 vccd2 _4906_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_62_94 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_62_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5886_ _5886_/A _5886_/B _5886_/C _5886_/D vssd2 vssd2 vccd2 vccd2 _5886_/X sky130_fd_sc_hd__or4_1
X_4837_ _4837_/A _4837_/B vssd2 vssd2 vccd2 vccd2 _4839_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_75_576 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_47_289 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7625_ _7627_/A vssd2 vssd2 vccd2 vccd2 _7625_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_105_317 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_90_568 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4768_ _4768_/A _4768_/B vssd2 vssd2 vccd2 vccd2 _4769_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_62_259 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7556_ _7557_/A vssd2 vssd2 vccd2 vccd2 _7556_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_153 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6507_ _6507_/A _6507_/B vssd2 vssd2 vccd2 vccd2 _6520_/A sky130_fd_sc_hd__xor2_2
X_4699_ _4699_/A _4699_/B vssd2 vssd2 vccd2 vccd2 _4700_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5009__D _5076_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_43_495 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7487_ _7524_/A vssd2 vssd2 vccd2 vccd2 _7487_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_164 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_113_361 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6438_ _6438_/A _6438_/B vssd2 vssd2 vccd2 vccd2 _6441_/A sky130_fd_sc_hd__xnor2_2
X_6369_ _6369_/A _6369_/B vssd2 vssd2 vccd2 vccd2 _6372_/A sky130_fd_sc_hd__xnor2_2
Xhold22 hold22/A vssd2 vssd2 vccd2 vccd2 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 hold11/A vssd2 vssd2 vccd2 vccd2 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6418__A _6855_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold33 hold33/A vssd2 vssd2 vccd2 vccd2 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd2 vssd2 vccd2 vccd2 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd2 vssd2 vccd2 vccd2 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd2 vssd2 vccd2 vccd2 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd2 vssd2 vccd2 vccd2 hold99/X sky130_fd_sc_hd__buf_1
Xhold88 hold88/A vssd2 vssd2 vccd2 vccd2 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd2 vssd2 vccd2 vccd2 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4661__A2 _5099_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4880__B _4880_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6153__A _6283_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_38_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_108_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_81_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_26_407 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_81_535 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_108_177 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__7115__B2 _7197_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_34_495 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA_8 hold73/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_21_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_21_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_318 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4120__B _5030_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_83_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_16_21 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_76_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_69_370 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5740_ _6282_/A _5755_/C _5739_/Y _6093_/A vssd2 vssd2 vccd2 vccd2 _5763_/B sky130_fd_sc_hd__a22o_1
XTAP_1090 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_576 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_57_565 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_8_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_72_557 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7410_ hold107/X _7674_/Q _7418_/S vssd2 vssd2 vccd2 vccd2 _7410_/X sky130_fd_sc_hd__mux2_1
X_5671_ _5811_/B _7855_/Q vssd2 vssd2 vccd2 vccd2 _5671_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_114_125 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_44_259 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4622_ _4622_/A _4622_/B vssd2 vssd2 vccd2 vccd2 _7738_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_309 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_52_270 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xmax_cap211 _4044_/B vssd2 vssd2 vccd2 vccd2 _4881_/A2 sky130_fd_sc_hd__buf_4
X_7341_ _7341_/A _7341_/B _7341_/C _7341_/D vssd2 vssd2 vccd2 vccd2 _7345_/A sky130_fd_sc_hd__or4_1
X_4553_ _4482_/A _4482_/B _4309_/B _4362_/B _4424_/A vssd2 vssd2 vccd2 vccd2 _4556_/B
+ sky130_fd_sc_hd__a2111o_2
XFILLER_0_40_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_114_169 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7272_ _7273_/A _7273_/B vssd2 vssd2 vccd2 vccd2 _7303_/B sky130_fd_sc_hd__nor2_1
Xhold536 la_data_in[31] vssd2 vssd2 vccd2 vccd2 hold55/A sky130_fd_sc_hd__dlygate4sd3_1
X_4484_ _4484_/A _4484_/B vssd2 vssd2 vccd2 vccd2 _7736_/D sky130_fd_sc_hd__xnor2_1
Xhold525 hold59/X vssd2 vssd2 vccd2 vccd2 input16/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 input19/X vssd2 vssd2 vccd2 vccd2 hold46/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold503 hold48/X vssd2 vssd2 vccd2 vccd2 _7866_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_454 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold547 hold70/X vssd2 vssd2 vccd2 vccd2 _7852_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 input24/X vssd2 vssd2 vccd2 vccd2 hold50/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 hold85/X vssd2 vssd2 vccd2 vccd2 input8/A sky130_fd_sc_hd__dlygate4sd3_1
X_6223_ _6100_/D _6587_/B _6222_/X _6220_/X _6281_/C vssd2 vssd2 vccd2 vccd2 _6223_/X
+ sky130_fd_sc_hd__a32o_2
XANTENNA__7622__A _7627_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4965__B _4965_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_852 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _6154_/A _6155_/B vssd2 vssd2 vccd2 vccd2 _6154_/Y sky130_fd_sc_hd__nor2_1
X_6085_ _6086_/A _6086_/B vssd2 vssd2 vccd2 vccd2 _6177_/A sky130_fd_sc_hd__and2_1
XFILLER_0_57_94 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_874 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4891__A2 _5315_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_863 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _5164_/A _5105_/B _5105_/C vssd2 vssd2 vccd2 vccd2 _5178_/B sky130_fd_sc_hd__nor3_2
XANTENNA__5142__A _5207_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5036_ _5035_/B _5035_/C _5035_/A vssd2 vssd2 vccd2 vccd2 _5037_/B sky130_fd_sc_hd__a21oi_1
XTAP_896 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout288_A _7629_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_32_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6987_ _7045_/A _7253_/A _6988_/A vssd2 vssd2 vccd2 vccd2 _7070_/A sky130_fd_sc_hd__or3_1
X_5938_ _6100_/D _6587_/B _5938_/C _5938_/D vssd2 vssd2 vccd2 vccd2 _5938_/X sky130_fd_sc_hd__and4_1
XANTENNA__6404__C _6404_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_90_321 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5869_ _7336_/A _5967_/A vssd2 vssd2 vccd2 vccd2 _5918_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_105_125 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_90_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_63_579 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7608_ _7613_/A vssd2 vssd2 vccd2 vccd2 _7608_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6553__C1 _5781_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7539_ _7561_/A vssd2 vssd2 vccd2 vccd2 _7539_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_495 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_105_169 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_31_421 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5317__A _5431_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7532__A _7564_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4331__A1 _4809_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_98_465 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_58_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_53_19 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_58_329 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_58_318 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XPHY_151 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_140 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_109_464 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_93_181 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_184 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_173 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_162 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6544__C1 _5736_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_26_259 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6330__B _6404_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_81_376 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_78_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_22_443 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_1_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7442__A _7452_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_94_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_27_64 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6910_ _7033_/A _7033_/C _7034_/A vssd2 vssd2 vccd2 vccd2 _6911_/B sky130_fd_sc_hd__a21oi_1
X_6841_ _6841_/A _6841_/B vssd2 vssd2 vccd2 vccd2 _6909_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_498 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_76_115 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_43_52 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_9_426 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_9_404 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4306__A _5548_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6772_ _6758_/A _6758_/B _6756_/X vssd2 vssd2 vccd2 vccd2 _6839_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_45_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3984_ _4214_/B _5030_/A _4162_/A _7775_/Q vssd2 vssd2 vccd2 vccd2 _3989_/D sky130_fd_sc_hd__and4b_1
XFILLER_0_45_535 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5723_ _5944_/B _5769_/B vssd2 vssd2 vccd2 vccd2 _5723_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_72_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5654_ _7847_/Q _7855_/Q _6019_/C vssd2 vssd2 vccd2 vccd2 _5655_/C sky130_fd_sc_hd__and3_1
XANTENNA__7336__B _7336_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4605_ _4605_/A _4605_/B vssd2 vssd2 vccd2 vccd2 _4606_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_32_218 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold311 hold664/X vssd2 vssd2 vccd2 vccd2 hold665/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold300 hold300/A vssd2 vssd2 vccd2 vccd2 la_data_out[16] sky130_fd_sc_hd__buf_12
X_7324_ _7324_/A _7324_/B vssd2 vssd2 vccd2 vccd2 _7334_/C sky130_fd_sc_hd__xor2_4
X_5585_ _5645_/B _5586_/B vssd2 vssd2 vccd2 vccd2 _6629_/C sky130_fd_sc_hd__and2_1
XFILLER_0_13_443 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4041__A _4454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_25_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_102_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4536_ _4393_/A _4393_/B _4468_/B _4469_/B _4469_/A vssd2 vssd2 vccd2 vccd2 _4538_/B
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout203_A _4217_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold333 _7746_/Q vssd2 vssd2 vccd2 vccd2 hold333/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold344 _7478_/X vssd2 vssd2 vccd2 vccd2 _7718_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold322 _7484_/X vssd2 vssd2 vccd2 vccd2 _7724_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_476 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_40_262 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4467_ _4467_/A _4467_/B vssd2 vssd2 vccd2 vccd2 _4468_/B sky130_fd_sc_hd__xnor2_2
X_7255_ _7291_/A _7255_/B vssd2 vssd2 vccd2 vccd2 _7256_/B sky130_fd_sc_hd__nor2_1
Xhold366 hold680/X vssd2 vssd2 vccd2 vccd2 _7780_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 _7653_/Q vssd2 vssd2 vccd2 vccd2 hold377/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 _7672_/Q vssd2 vssd2 vccd2 vccd2 hold355/X sky130_fd_sc_hd__dlygate4sd3_1
X_6206_ _6206_/A _6206_/B vssd2 vssd2 vccd2 vccd2 _6208_/B sky130_fd_sc_hd__xnor2_2
X_7186_ _7186_/A _7186_/B vssd2 vssd2 vccd2 vccd2 _7188_/B sky130_fd_sc_hd__xnor2_1
X_4398_ _5029_/A _4966_/A vssd2 vssd2 vccd2 vccd2 _4401_/A sky130_fd_sc_hd__or2_2
Xhold388 _7675_/Q vssd2 vssd2 vccd2 vccd2 hold388/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 _7682_/Q vssd2 vssd2 vccd2 vccd2 hold399/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4313__A1 _7766_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6137_ _5778_/X _5786_/Y _6973_/B _5736_/X vssd2 vssd2 vccd2 vccd2 _6139_/A sky130_fd_sc_hd__a211o_1
XTAP_660 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _6068_/A _6068_/B _6067_/A vssd2 vssd2 vccd2 vccd2 _6189_/A sky130_fd_sc_hd__or3b_2
XANTENNA__5813__A1 _7844_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5019_ _5021_/A _5021_/B vssd2 vssd2 vccd2 vccd2 _5019_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_95_424 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4861__D _5076_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_48_362 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5041__A2 _5374_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_36_546 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_63_332 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__7527__A _7563_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_36_579 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_63_387 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_51_516 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_467 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_90_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6150__B _6150_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_16_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_101_161 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_64_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5804__A1 _7847_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_98_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_59_627 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_86_435 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6044__C _6939_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_67_671 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_58_159 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_13_11 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_362 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_66_181 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6780__A2 _7222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_109_261 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6341__A _6855_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_89_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_54_343 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_42_516 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_42_549 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5370_ _5370_/A _5370_/B _5370_/C vssd2 vssd2 vccd2 vccd2 _5371_/B sky130_fd_sc_hd__or3_1
XANTENNA__4796__A _5029_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4321_ _4367_/B _4321_/B vssd2 vssd2 vccd2 vccd2 _4323_/C sky130_fd_sc_hd__and2_1
XFILLER_0_22_295 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7040_ _7040_/A _7040_/B vssd2 vssd2 vccd2 vccd2 _7042_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_10_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4252_ _4490_/A _4252_/B _4252_/C _4252_/D vssd2 vssd2 vccd2 vccd2 _4252_/X sky130_fd_sc_hd__or4_1
XANTENNA__5404__B _5498_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4183_ _4183_/A _4183_/B vssd2 vssd2 vccd2 vccd2 _4186_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_77_413 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4962__C _5406_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_77_457 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_77_446 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7873_ _7878_/CLK _7873_/D _7632_/Y vssd2 vssd2 vccd2 vccd2 _7873_/Q sky130_fd_sc_hd__dfrtp_2
X_6824_ _6825_/A _6825_/B vssd2 vssd2 vccd2 vccd2 _6824_/X sky130_fd_sc_hd__or2_1
XANTENNA__6220__A1 _6093_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_92_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6755_ _6689_/A _6689_/B _6687_/Y vssd2 vssd2 vccd2 vccd2 _6757_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_9_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3967_ _4018_/A _4018_/B _3967_/C _3967_/D vssd2 vssd2 vccd2 vccd2 _3967_/X sky130_fd_sc_hd__and4b_1
XANTENNA__6220__B2 _6253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6251__A _6402_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_45_343 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5706_ _6510_/B _6670_/B vssd2 vssd2 vccd2 vccd2 _5850_/B sky130_fd_sc_hd__nor2_2
X_6686_ _6604_/A _6604_/B _6602_/X vssd2 vssd2 vccd2 vccd2 _6688_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_5_440 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3898_ _4326_/D _4002_/B _3898_/C vssd2 vssd2 vccd2 vccd2 _3898_/X sky130_fd_sc_hd__and3_1
XFILLER_0_33_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_60_357 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5637_ _5638_/B _5638_/C vssd2 vssd2 vccd2 vccd2 _5661_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_484 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5568_ _5553_/A _5553_/B _5567_/X vssd2 vssd2 vccd2 vccd2 _5568_/Y sky130_fd_sc_hd__a21boi_1
X_7307_ _7309_/A vssd2 vssd2 vccd2 vccd2 _7307_/Y sky130_fd_sc_hd__inv_2
Xhold130 hold387/X vssd2 vssd2 vccd2 vccd2 _7769_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 wbs_dat_i[0] vssd2 vssd2 vccd2 vccd2 input83/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 hold357/X vssd2 vssd2 vccd2 vccd2 _7799_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4519_ _4656_/A _4519_/B _4519_/C vssd2 vssd2 vccd2 vccd2 _4519_/X sky130_fd_sc_hd__and3_1
XANTENNA__7082__A _7082_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7238_ _7239_/B _7239_/C _7239_/A vssd2 vssd2 vccd2 vccd2 _7270_/A sky130_fd_sc_hd__o21ai_1
Xhold163 _7445_/X vssd2 vssd2 vccd2 vccd2 _7446_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7484__B1 _7485_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold174 wbs_dat_i[1] vssd2 vssd2 vccd2 vccd2 input90/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _7363_/X vssd2 vssd2 vccd2 vccd2 _7364_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ _5499_/A _5499_/B vssd2 vssd2 vccd2 vccd2 _5500_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_111_492 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold196 hold395/X vssd2 vssd2 vccd2 vccd2 _7795_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7169_ _7169_/A _7169_/B _7169_/C vssd2 vssd2 vccd2 vccd2 _7214_/B sky130_fd_sc_hd__nand3_2
XTAP_490 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6039__B2 _6093_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1623 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6145__B _6738_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4591__D _5222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_83_416 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_48_170 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_63_151 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_253 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_59_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7475__B1 _7483_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_91_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4782__C _5099_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_435 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_59_424 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_10 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_24_21 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_86_265 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_86_243 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_4870_ _4966_/A _5276_/A _4781_/X _4783_/B vssd2 vssd2 vccd2 vccd2 _4872_/B sky130_fd_sc_hd__o31a_1
X_3821_ _3821_/A _7804_/Q vssd2 vssd2 vccd2 vccd2 _3821_/X sky130_fd_sc_hd__or2_1
X_6540_ _6489_/A _6489_/B _6490_/X vssd2 vssd2 vccd2 vccd2 _6542_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_490 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__6071__A _6670_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_42_313 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_15_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_15_516 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_387 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6471_ _6422_/A _6422_/B _6420_/Y vssd2 vssd2 vccd2 vccd2 _6489_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_2_410 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5422_ _5472_/A _5422_/B _5465_/A vssd2 vssd2 vccd2 vccd2 _5424_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_112_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5353_ _5353_/A _5353_/B vssd2 vssd2 vccd2 vccd2 _5445_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_112_289 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4304_ _4304_/A _4304_/B vssd2 vssd2 vccd2 vccd2 _4308_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__7466__B1 _7485_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5284_ _5284_/A _5341_/A vssd2 vssd2 vccd2 vccd2 _5287_/A sky130_fd_sc_hd__or2_1
X_7023_ _7023_/A vssd2 vssd2 vccd2 vccd2 _7083_/A sky130_fd_sc_hd__inv_2
X_4235_ _4237_/A _4237_/B vssd2 vssd2 vccd2 vccd2 _4235_/X sky130_fd_sc_hd__and2_1
XANTENNA__7630__A _7641_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4166_ _4162_/X _4165_/Y _4057_/C vssd2 vssd2 vccd2 vccd2 _4166_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5150__A _5276_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4097_ _5455_/A _4193_/A vssd2 vssd2 vccd2 vccd2 _4139_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4894__A2_N _5550_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_77_243 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7856_ _7886_/CLK _7856_/D _7615_/Y vssd2 vssd2 vccd2 vccd2 _7856_/Q sky130_fd_sc_hd__dfrtp_4
X_6807_ _6876_/B _6806_/C _6806_/A vssd2 vssd2 vccd2 vccd2 _6808_/C sky130_fd_sc_hd__a21o_1
X_7787_ _7787_/CLK _7787_/D _7546_/Y vssd2 vssd2 vccd2 vccd2 _7787_/Q sky130_fd_sc_hd__dfrtp_2
X_4999_ _5133_/A _4999_/B vssd2 vssd2 vccd2 vccd2 _7743_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_321 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6738_ _6738_/A _7099_/B vssd2 vssd2 vccd2 vccd2 _6739_/B sky130_fd_sc_hd__nand2_1
X_6669_ _6670_/A _6670_/B vssd2 vssd2 vccd2 vccd2 _6669_/X sky130_fd_sc_hd__and2_4
XFILLER_0_45_173 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7457__B1 _7485_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6432__A1 _6093_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1431 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_265 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5210__D _5498_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1475 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3946__C _7768_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_36_151 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_24_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_10_45 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_17_wb_clk_i clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7768_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7160__A2 _7255_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4777__C _5142_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_20_530 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_20_563 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4496__D _4782_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_19_32 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_19_43 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7450__A _7450_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4020_ _4214_/C _4020_/B _4122_/D vssd2 vssd2 vccd2 vccd2 _4020_/X sky130_fd_sc_hd__and3_1
X_5971_ _7336_/A _5968_/A _5968_/X _6011_/A vssd2 vssd2 vccd2 vccd2 _7811_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_35_64 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4922_ _4923_/A _4923_/B _4923_/C vssd2 vssd2 vccd2 vccd2 _4922_/X sky130_fd_sc_hd__a21o_1
X_7710_ _7771_/CLK _7710_/D vssd2 vssd2 vccd2 vccd2 _7710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_596 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_74_202 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7641_ _7641_/A vssd2 vssd2 vccd2 vccd2 _7641_/Y sky130_fd_sc_hd__inv_2
X_4853_ _4854_/A _4854_/B _4854_/C vssd2 vssd2 vccd2 vccd2 _4990_/A sky130_fd_sc_hd__o21a_2
XANTENNA__6187__B1 _6069_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_74_235 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6513__B _7294_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_51_52 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_7_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7572_ _7613_/A vssd2 vssd2 vccd2 vccd2 _7572_/Y sky130_fd_sc_hd__inv_2
X_4784_ _4966_/A _5276_/A vssd2 vssd2 vccd2 vccd2 _4785_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_27_151 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_28_674 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3804_ _3804_/A vssd2 vssd2 vccd2 vccd2 _5586_/B sky130_fd_sc_hd__clkinv_4
X_6523_ _6523_/A _6523_/B vssd2 vssd2 vccd2 vccd2 _6524_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_55_482 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_15_313 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_27_173 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6454_ _6455_/A _6455_/B vssd2 vssd2 vccd2 vccd2 _6537_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_15_368 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7625__A _7627_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_70_485 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_30_327 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5405_ _5403_/X _5405_/B vssd2 vssd2 vccd2 vccd2 _5407_/A sky130_fd_sc_hd__and2b_1
X_6385_ _6387_/C vssd2 vssd2 vccd2 vccd2 _6385_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_62_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__5145__A _5145_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_11_552 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_23_390 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_30_349 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5336_ _5336_/A _5336_/B vssd2 vssd2 vccd2 vccd2 _5339_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_11_574 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_76_60 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5267_ _5267_/A _5267_/B vssd2 vssd2 vccd2 vccd2 _5270_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7006_ _7007_/A _7007_/B _7007_/C vssd2 vssd2 vccd2 vccd2 _7012_/A sky130_fd_sc_hd__a21oi_1
X_4218_ _4598_/A _4662_/B _4219_/B vssd2 vssd2 vccd2 vccd2 _4220_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__7360__A _7436_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5907__A_N _6138_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5198_ _5198_/A _5357_/B vssd2 vssd2 vccd2 vccd2 _7746_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_305 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4149_ _4149_/A _4149_/B _4149_/C vssd2 vssd2 vccd2 vccd2 _4149_/X sky130_fd_sc_hd__or3_1
XANTENNA__4208__B _4966_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_93_533 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_93_500 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_38_427 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6423__B _7094_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7839_ _7870_/CLK _7839_/D _7598_/Y vssd2 vssd2 vccd2 vccd2 _7839_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_73_290 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_33_121 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7535__A _7557_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_33_154 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_104_554 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__7142__A2 _7294_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_104_598 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_104_587 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5205__D _5498_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout292 _7629_/A vssd2 vssd2 vccd2 vccd2 _7613_/A sky130_fd_sc_hd__buf_6
Xfanout281 _7557_/A vssd2 vssd2 vccd2 vccd2 _7524_/A sky130_fd_sc_hd__buf_8
Xfanout270 _7773_/Q vssd2 vssd2 vccd2 vccd2 _4656_/A sky130_fd_sc_hd__buf_4
XTAP_1250 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3957__B _5030_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_29_438 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1272 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_533 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_29_449 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1294 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_216 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_4_527 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_97_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_52_474 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_40_625 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_110_557 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6170_ _6111_/A _6111_/C _6111_/B vssd2 vssd2 vccd2 vccd2 _6172_/B sky130_fd_sc_hd__a21bo_1
X_5121_ _5122_/A _5122_/B vssd2 vssd2 vccd2 vccd2 _5121_/X sky130_fd_sc_hd__or2_1
XANTENNA__6508__B _7099_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5052_ _5052_/A _5052_/B vssd2 vssd2 vccd2 vccd2 _5055_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_46_41 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4309__A _5455_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4003_ _4656_/B _5458_/A _4100_/B vssd2 vssd2 vccd2 vccd2 _4004_/B sky130_fd_sc_hd__and3_1
XANTENNA__6227__C _7197_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_75_522 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5954_ _6402_/A _6150_/A _5909_/A _5908_/A vssd2 vssd2 vccd2 vccd2 _5956_/C sky130_fd_sc_hd__a31oi_2
XANTENNA__5080__B1 _5468_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_4905_ _4822_/A _4822_/B _4820_/Y vssd2 vssd2 vccd2 vccd2 _4907_/B sky130_fd_sc_hd__o21ba_2
X_5885_ _6074_/A _5977_/B _5884_/X vssd2 vssd2 vccd2 vccd2 _5885_/X sky130_fd_sc_hd__a21o_1
X_4836_ _4837_/A _4837_/B vssd2 vssd2 vccd2 vccd2 _4923_/A sky130_fd_sc_hd__or2_1
XFILLER_0_75_588 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_47_257 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_28_460 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4044__A _4044_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7624_ _7627_/A vssd2 vssd2 vccd2 vccd2 _7624_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_62_249 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_15_110 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7555_ _7563_/A vssd2 vssd2 vccd2 vccd2 _7555_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_105_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6506_ _6581_/A _7045_/A vssd2 vssd2 vccd2 vccd2 _6507_/B sky130_fd_sc_hd__nor2_1
X_4767_ _4767_/A _4767_/B vssd2 vssd2 vccd2 vccd2 _4768_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_43_430 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_15_121 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4698_ _4699_/A _4699_/B vssd2 vssd2 vccd2 vccd2 _4839_/A sky130_fd_sc_hd__or2_1
XFILLER_0_43_485 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7486_ _7726_/Q _7453_/Y hold104/X hold697/X vssd2 vssd2 vccd2 vccd2 _7486_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_113_373 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6437_ _6437_/A _6437_/B vssd2 vssd2 vccd2 vccd2 _6438_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_293 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6368_ _6368_/A _6368_/B vssd2 vssd2 vccd2 vccd2 _6369_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_87_81 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5319_ _5320_/A _5320_/B vssd2 vssd2 vccd2 vccd2 _5370_/B sky130_fd_sc_hd__and2_1
X_6299_ _6299_/A _6299_/B vssd2 vssd2 vccd2 vccd2 _6302_/A sky130_fd_sc_hd__xnor2_2
Xhold23 hold23/A vssd2 vssd2 vccd2 vccd2 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 hold12/A vssd2 vssd2 vccd2 vccd2 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6418__B _7037_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold34 hold34/A vssd2 vssd2 vccd2 vccd2 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd2 vssd2 vccd2 vccd2 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd2 vssd2 vccd2 vccd2 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd2 vssd2 vccd2 vccd2 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd2 vssd2 vccd2 vccd2 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd2 vssd2 vccd2 vccd2 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4219__A _4598_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_113 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_66_511 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_78_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_66_555 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_66_533 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6153__B _6281_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_38_235 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_66_577 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_19_460 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_26_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_38_257 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_81_558 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_81_547 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5992__B _5992_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_108_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__3793__A _4656_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_9 la_data_in[3] vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_21_146 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6874__A1 _6738_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_319 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_614 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_83_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_107_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_88_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_88_146 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_69_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_72_503 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1091 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_588 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_17_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5670_ _5811_/B _5811_/C _5878_/B _5669_/X vssd2 vssd2 vccd2 vccd2 _5670_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_29_257 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_84_396 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_72_525 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4621_ _4621_/A _4621_/B vssd2 vssd2 vccd2 vccd2 _4622_/B sky130_fd_sc_hd__and2_1
XFILLER_0_25_441 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_114_137 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7340_ _7340_/A _7340_/B _7340_/C _7340_/D vssd2 vssd2 vccd2 vccd2 _7340_/X sky130_fd_sc_hd__or4_1
X_4552_ _4619_/B _4552_/B vssd2 vssd2 vccd2 vccd2 _4556_/A sky130_fd_sc_hd__and2_2
X_7271_ _7303_/A _7271_/B vssd2 vssd2 vccd2 vccd2 _7273_/B sky130_fd_sc_hd__or2_1
Xmax_cap234 _5921_/D vssd2 vssd2 vccd2 vccd2 _6019_/D sky130_fd_sc_hd__buf_2
X_4483_ _5455_/A _4424_/A _4424_/B vssd2 vssd2 vccd2 vccd2 _4484_/B sky130_fd_sc_hd__a21oi_1
Xhold504 la_data_in[11] vssd2 vssd2 vccd2 vccd2 hold11/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold526 input16/X vssd2 vssd2 vccd2 vccd2 hold60/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 hold46/X vssd2 vssd2 vccd2 vccd2 _7865_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_433 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_40_444 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_110_321 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold537 hold55/X vssd2 vssd2 vccd2 vccd2 input25/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 hold50/X vssd2 vssd2 vccd2 vccd2 _7869_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 la_data_in[22] vssd2 vssd2 vccd2 vccd2 hold71/A sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap245 _4068_/B vssd2 vssd2 vccd2 vccd2 _4815_/B sky130_fd_sc_hd__buf_6
X_6222_ _6510_/A _5937_/B _5938_/C _6094_/B _6283_/A vssd2 vssd2 vccd2 vccd2 _6222_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_110_365 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_853 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _6283_/A _6281_/B _6281_/C vssd2 vssd2 vccd2 vccd2 _6153_/X sky130_fd_sc_hd__and3_2
X_6084_ _6144_/A _6084_/B vssd2 vssd2 vccd2 vccd2 _6086_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_57_84 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_875 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _5104_/A _5104_/B vssd2 vssd2 vccd2 vccd2 _5105_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__5142__B _5431_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5035_ _5035_/A _5035_/B _5035_/C vssd2 vssd2 vccd2 vccd2 _5091_/B sky130_fd_sc_hd__and3_1
XTAP_897 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout183_A _6103_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_79_124 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_79_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__3878__A _4454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_95_617 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_79_179 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6986_ _6986_/A _7253_/A vssd2 vssd2 vccd2 vccd2 _6988_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_87_190 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_75_330 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5937_ _6157_/A _5937_/B vssd2 vssd2 vccd2 vccd2 _5938_/D sky130_fd_sc_hd__and2_1
XANTENNA__6404__D _6404_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_63_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_90_333 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5868_ _7807_/D _5868_/B _5868_/C vssd2 vssd2 vccd2 vccd2 _5967_/A sky130_fd_sc_hd__or3_1
XFILLER_0_63_525 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7607_ _7613_/A vssd2 vssd2 vccd2 vccd2 _7607_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_35_216 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_638 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4819_ _4819_/A _4819_/B vssd2 vssd2 vccd2 vccd2 _4821_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__6553__B1 _7143_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_16_441 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5799_ _6253_/B _6253_/C _6018_/D _5811_/B vssd2 vssd2 vccd2 vccd2 _5977_/B sky130_fd_sc_hd__and4_2
XFILLER_0_105_137 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_43_260 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7538_ _7557_/A vssd2 vssd2 vccd2 vccd2 _7538_/Y sky130_fd_sc_hd__inv_2
X_7469_ _7709_/Q _7483_/A2 _7483_/B1 hold325/X vssd2 vssd2 vccd2 vccd2 _7469_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_31_433 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5317__B _5550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_113_181 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_3_390 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_31_499 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_98_400 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_85_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_1_1__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_85_127 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_152 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_130 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_185 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_174 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_163 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_54_547 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_54_525 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_26_227 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_196 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_93_193 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6544__B1 _7253_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_105_671 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_1_349 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_22_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_94_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_89_466 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6840_ _6768_/A _6768_/B _6762_/A vssd2 vssd2 vccd2 vccd2 _6841_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_43_20 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6771_ _6909_/A _6771_/B vssd2 vssd2 vccd2 vccd2 _7823_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_149 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_9_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3983_ _4214_/C _4164_/C vssd2 vssd2 vccd2 vccd2 _3989_/C sky130_fd_sc_hd__nor2_1
X_5722_ _6152_/B _5937_/B vssd2 vssd2 vccd2 vccd2 _5944_/D sky130_fd_sc_hd__nor2_1
XANTENNA__6802__A _6973_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_5_611 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5653_ _7843_/Q _7855_/Q _5653_/C _6016_/B vssd2 vssd2 vccd2 vccd2 _5653_/X sky130_fd_sc_hd__and4_1
X_4604_ _4605_/A _4605_/B vssd2 vssd2 vccd2 vccd2 _4604_/X sky130_fd_sc_hd__and2_1
X_5584_ _5583_/A _5583_/B _5645_/B vssd2 vssd2 vccd2 vccd2 _5584_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_0_5_644 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold301 hold654/X vssd2 vssd2 vccd2 vccd2 hold655/A sky130_fd_sc_hd__dlygate4sd3_1
X_7323_ _7324_/A _7324_/B vssd2 vssd2 vccd2 vccd2 _7334_/B sky130_fd_sc_hd__nand2b_1
X_4535_ _4535_/A _4535_/B vssd2 vssd2 vccd2 vccd2 _4538_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_591 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xhold312 hold312/A vssd2 vssd2 vccd2 vccd2 la_data_out[25] sky130_fd_sc_hd__buf_12
Xhold334 _7474_/X vssd2 vssd2 vccd2 vccd2 _7714_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _7740_/Q vssd2 vssd2 vccd2 vccd2 hold323/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7633__A _7641_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_40_230 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_68_50 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4466_ _4467_/A _4467_/B vssd2 vssd2 vccd2 vccd2 _4534_/A sky130_fd_sc_hd__and2b_1
X_7254_ _7252_/X _7254_/B vssd2 vssd2 vccd2 vccd2 _7256_/A sky130_fd_sc_hd__and2b_1
Xhold345 _7753_/Q vssd2 vssd2 vccd2 vccd2 hold345/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 hold690/X vssd2 vssd2 vccd2 vccd2 _7759_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_488 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold367 _7656_/Q vssd2 vssd2 vccd2 vccd2 hold367/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 _7693_/Q vssd2 vssd2 vccd2 vccd2 hold356/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_285 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6205_ _6634_/B _6571_/A vssd2 vssd2 vccd2 vccd2 _6206_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_68_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7185_ _7186_/B _7186_/A vssd2 vssd2 vccd2 vccd2 _7232_/A sky130_fd_sc_hd__nand2b_1
X_4397_ _4896_/A _5030_/B _5030_/A vssd2 vssd2 vccd2 vccd2 _4402_/A sky130_fd_sc_hd__and3b_2
Xhold389 _7694_/Q vssd2 vssd2 vccd2 vccd2 hold389/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6136_ _6550_/A _7037_/A vssd2 vssd2 vccd2 vccd2 _6140_/A sky130_fd_sc_hd__nor2_1
XTAP_650 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _6067_/A _6067_/B vssd2 vssd2 vccd2 vccd2 _7813_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__4077__B2 _4328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5018_ _4941_/A _4943_/B _4941_/B vssd2 vssd2 vccd2 vccd2 _5021_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_95_436 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_67_127 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6969_ _7025_/D _6969_/B vssd2 vssd2 vccd2 vccd2 _7033_/D sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_352 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_75_182 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_402 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4001__A1 _7761_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5328__A _5328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4001__B2 _7762_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_606 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6044__D _6989_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_13_23 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_39_374 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_109_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6341__B _6973_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_66_193 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_89_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_50_550 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5740__A1 _6282_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5740__B2 _6093_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_1_124 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4796__B _5406_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4320_ _4598_/A _4782_/B _4319_/B vssd2 vssd2 vccd2 vccd2 _4321_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_425 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_10_414 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6069__A _6069_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4251_ _4656_/A _4251_/B vssd2 vssd2 vccd2 vccd2 _4251_/X sky130_fd_sc_hd__and2_1
XANTENNA__5404__C _5468_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4182_ _4183_/A _4183_/B vssd2 vssd2 vccd2 vccd2 _4237_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_38_75 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4059__B2 _7767_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_54_41 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7872_ _7878_/CLK _7872_/D _7631_/Y vssd2 vssd2 vccd2 vccd2 _7872_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5008__B1 _5076_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_54_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6823_ _6746_/A _6746_/B _6744_/X vssd2 vssd2 vccd2 vccd2 _6825_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__7628__A _7629_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6754_ _6754_/A _6754_/B vssd2 vssd2 vccd2 vccd2 _6757_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3966_ _7772_/Q _3965_/A _3965_/Y _4809_/A vssd2 vssd2 vccd2 vccd2 _3967_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_18_514 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6220__A2 _6281_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6251__B _7143_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6685_ _6685_/A _6685_/B vssd2 vssd2 vccd2 vccd2 _6688_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_193 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5705_ _7885_/Q _5694_/X _5705_/C _5735_/B vssd2 vssd2 vccd2 vccd2 _6670_/B sky130_fd_sc_hd__and4bb_4
XFILLER_0_18_569 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_92_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_72_163 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_72_141 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_60_314 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5636_ _5638_/B _5638_/C vssd2 vssd2 vccd2 vccd2 _5811_/C sky130_fd_sc_hd__and2_2
X_3897_ _7791_/Q _4328_/A _4148_/B _4080_/D vssd2 vssd2 vccd2 vccd2 _3898_/C sky130_fd_sc_hd__and4_1
XFILLER_0_33_517 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5567_ _5458_/A _5431_/B _5550_/B _4814_/B _5529_/B vssd2 vssd2 vccd2 vccd2 _5567_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_82 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7306_ _7306_/A _7306_/B vssd2 vssd2 vccd2 vccd2 _7309_/A sky130_fd_sc_hd__nor2_1
X_4518_ _4736_/A _5220_/A vssd2 vssd2 vccd2 vccd2 _4532_/A sky130_fd_sc_hd__or2_1
Xhold131 _7373_/X vssd2 vssd2 vccd2 vccd2 _7374_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 _7437_/X vssd2 vssd2 vccd2 vccd2 _7438_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 input83/X vssd2 vssd2 vccd2 vccd2 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 wbs_dat_i[8] vssd2 vssd2 vccd2 vccd2 input97/A sky130_fd_sc_hd__dlygate4sd3_1
X_5498_ _5498_/A _5550_/A _5528_/A _5498_/D vssd2 vssd2 vccd2 vccd2 _5499_/B sky130_fd_sc_hd__or4_1
XANTENNA__7082__B _7082_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7237_ _7237_/A _7291_/B vssd2 vssd2 vccd2 vccd2 _7239_/C sky130_fd_sc_hd__nor2_1
X_4449_ _4449_/A _4449_/B vssd2 vssd2 vccd2 vccd2 _4451_/B sky130_fd_sc_hd__xnor2_4
Xhold186 wbs_dat_i[2] vssd2 vssd2 vccd2 vccd2 input91/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 input90/X vssd2 vssd2 vccd2 vccd2 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 hold361/X vssd2 vssd2 vccd2 vccd2 _7791_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 _7429_/X vssd2 vssd2 vccd2 vccd2 _7430_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_81 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7168_ _7168_/A _7168_/B vssd2 vssd2 vccd2 vccd2 _7169_/C sky130_fd_sc_hd__xnor2_1
X_6119_ _6119_/A _6119_/B _6119_/C vssd2 vssd2 vccd2 vccd2 _6128_/B sky130_fd_sc_hd__or3_1
XANTENNA__6707__A _6707_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7099_ _7145_/A _7099_/B vssd2 vssd2 vccd2 vccd2 _7100_/B sky130_fd_sc_hd__nand2_1
XTAP_491 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6426__B _6426_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1624 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_428 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7538__A _7557_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_48_182 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_36_322 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_36_333 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_106_221 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_106_265 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_63_174 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_51_358 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_32_572 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_99_561 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_91_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4782__D _4965_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_99_583 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_24_33 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_24_44 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6352__A _6425_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_277 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7448__A _7450_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4213__A1 _4656_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3820_ _4745_/A _4522_/C vssd2 vssd2 vccd2 vccd2 _3820_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4213__B2 _4454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6470_ _5819_/B _7222_/A _6410_/B _6408_/X vssd2 vssd2 vccd2 vccd2 _6491_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_40_65 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6910__B1 _7034_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5421_ _5421_/A _5421_/B vssd2 vssd2 vccd2 vccd2 _5465_/A sky130_fd_sc_hd__or2_1
X_5352_ _5353_/B _5353_/A vssd2 vssd2 vccd2 vccd2 _5352_/X sky130_fd_sc_hd__and2b_1
XANTENNA__4600__A _4708_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_49_30 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_50_391 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_10_222 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4303_ _4303_/A _4303_/B _4303_/C _4303_/D vssd2 vssd2 vccd2 vccd2 _4360_/B sky130_fd_sc_hd__or4_1
X_7022_ _7024_/A _7024_/B vssd2 vssd2 vccd2 vccd2 _7023_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_74 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5283_ _5431_/A _5404_/A _5406_/A _5498_/A vssd2 vssd2 vccd2 vccd2 _5341_/A sky130_fd_sc_hd__nor4_2
X_4234_ _4234_/A _4234_/B vssd2 vssd2 vccd2 vccd2 _4237_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4165_ _4163_/Y _4164_/X _3986_/A vssd2 vssd2 vccd2 vccd2 _4165_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_65_62 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5431__A _5431_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5150__B _5414_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4096_ _4096_/A _4096_/B vssd2 vssd2 vccd2 vccd2 _4193_/A sky130_fd_sc_hd__or2_1
XANTENNA_fanout263_A _7850_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7855_ _7886_/CLK _7855_/D _7614_/Y vssd2 vssd2 vccd2 vccd2 _7855_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_288 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6806_ _6806_/A _6876_/B _6806_/C vssd2 vssd2 vccd2 vccd2 _6808_/B sky130_fd_sc_hd__nand3_1
XANTENNA__7358__A _7436_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_37_108 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4998_ _5548_/A _5133_/B vssd2 vssd2 vccd2 vccd2 _4999_/B sky130_fd_sc_hd__nor2_1
X_7786_ _7802_/CLK _7786_/D _7545_/Y vssd2 vssd2 vccd2 vccd2 _7786_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_61_601 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6737_ _6737_/A _6737_/B vssd2 vssd2 vccd2 vccd2 _6739_/A sky130_fd_sc_hd__nor2_1
X_3949_ _7776_/Q _7775_/Q _7777_/Q _4050_/B vssd2 vssd2 vccd2 vccd2 _3950_/B sky130_fd_sc_hd__o31a_2
X_6668_ _6668_/A _7294_/C vssd2 vssd2 vccd2 vccd2 _6673_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_325 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6599_ _6599_/A _6599_/B vssd2 vssd2 vccd2 vccd2 _6600_/B sky130_fd_sc_hd__xnor2_2
X_5619_ _7863_/Q _5619_/B vssd2 vssd2 vccd2 vccd2 _6075_/C sky130_fd_sc_hd__xor2_4
XANTENNA__4510__A _5029_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_60_188 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_60_177 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5325__B _5498_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_41_380 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_88_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4443__A1 _4810_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1432 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_119 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__3796__A _4162_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1498 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6735__A3 _7294_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_71_409 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_36_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_36_163 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_107_541 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_101_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_52_645 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_24_369 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4777__D _5076_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_20_553 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6671__A2 _7313_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5970_ _7336_/A _6068_/A vssd2 vssd2 vccd2 vccd2 _6011_/A sky130_fd_sc_hd__and2_1
XFILLER_0_59_222 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_59_200 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_35_54 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4921_ _4923_/A _4923_/B _4923_/C vssd2 vssd2 vccd2 vccd2 _4924_/A sky130_fd_sc_hd__a21oi_1
X_4852_ _4778_/A _4780_/B _4778_/B vssd2 vssd2 vccd2 vccd2 _4854_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__7178__A _7237_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7640_ _7641_/A vssd2 vssd2 vccd2 vccd2 _7640_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_74_247 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_3803_ _7842_/Q vssd2 vssd2 vccd2 vccd2 _3803_/Y sky130_fd_sc_hd__inv_2
X_7571_ _7613_/A vssd2 vssd2 vccd2 vccd2 _7571_/Y sky130_fd_sc_hd__inv_2
X_4783_ _4781_/X _4783_/B vssd2 vssd2 vccd2 vccd2 _4785_/A sky130_fd_sc_hd__and2b_1
X_6522_ _6523_/A _6523_/B vssd2 vssd2 vccd2 vccd2 _6522_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_55_494 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6453_ _6453_/A _6453_/B vssd2 vssd2 vccd2 vccd2 _6455_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_15_347 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_70_497 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_70_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5404_ _5404_/A _5498_/A _5468_/A _5498_/D vssd2 vssd2 vccd2 vccd2 _5405_/B sky130_fd_sc_hd__or4_1
XFILLER_0_42_188 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6384_ _6384_/A _6384_/B vssd2 vssd2 vccd2 vccd2 _6387_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__5145__B _5145_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_11_542 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_11_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5335_ _5379_/B _5335_/B vssd2 vssd2 vccd2 vccd2 _5336_/B sky130_fd_sc_hd__xor2_2
XANTENNA__7641__A _7641_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5266_ _5266_/A _5266_/B vssd2 vssd2 vccd2 vccd2 _5267_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__6257__A _6550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_76_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7005_ _7005_/A _7005_/B vssd2 vssd2 vccd2 vccd2 _7007_/C sky130_fd_sc_hd__xnor2_1
X_4217_ _4212_/X _4213_/X _4216_/X _4164_/C vssd2 vssd2 vccd2 vccd2 _4217_/Y sky130_fd_sc_hd__o31ai_4
X_5197_ _5250_/D _5197_/B vssd2 vssd2 vccd2 vccd2 _5357_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_97_317 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6634__A_N _6707_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4148_ _4457_/A _4148_/B _4148_/C _4148_/D vssd2 vssd2 vccd2 vccd2 _4148_/X sky130_fd_sc_hd__or4_1
XFILLER_0_78_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4079_ _4075_/X _4077_/X _4078_/X _4083_/B vssd2 vssd2 vccd2 vccd2 _4088_/A sky130_fd_sc_hd__o31ai_4
XFILLER_0_78_542 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7838_ _7838_/CLK _7838_/D _7597_/Y vssd2 vssd2 vccd2 vccd2 _7838_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_545 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_65_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_38_439 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_46_461 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7769_ _7802_/CLK _7769_/D _7528_/Y vssd2 vssd2 vccd2 vccd2 _7769_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__7127__B1 _7082_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_18_174 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_18_185 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_100 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_61_464 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_61_431 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_104_533 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_33_166 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_177 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6638__C1 _5781_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7551__A _7557_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout260 _7852_/Q vssd2 vssd2 vccd2 vccd2 _6397_/A sky130_fd_sc_hd__buf_2
Xfanout282 _7563_/A vssd2 vssd2 vccd2 vccd2 _7557_/A sky130_fd_sc_hd__buf_8
Xfanout271 _7773_/Q vssd2 vssd2 vccd2 vccd2 _4706_/A1 sky130_fd_sc_hd__buf_2
Xfanout293 input49/X vssd2 vssd2 vccd2 vccd2 _7629_/A sky130_fd_sc_hd__buf_8
XANTENNA__5613__B1 _5645_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1240 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_394 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1273 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_545 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1251 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_236 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1295 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_56_269 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_37_461 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_21_23 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_64_291 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_52_431 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_97_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_20_361 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_110_569 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5120_ _5060_/A _5060_/B _5058_/Y vssd2 vssd2 vccd2 vccd2 _5122_/B sky130_fd_sc_hd__a21oi_2
X_5051_ _5051_/A _5051_/B vssd2 vssd2 vccd2 vccd2 _5052_/B sky130_fd_sc_hd__xor2_4
X_4002_ _4002_/A _4002_/B _4002_/C vssd2 vssd2 vccd2 vccd2 _4002_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_94_309 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7400__S _7418_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5953_ _5952_/B _5952_/C _5952_/A vssd2 vssd2 vccd2 vccd2 _5956_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__5080__A1 _5210_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5080__B2 _5210_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_62_41 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_47_203 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_75_556 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_62_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4904_ _4904_/A _4904_/B vssd2 vssd2 vccd2 vccd2 _4907_/A sky130_fd_sc_hd__xnor2_4
X_5884_ _6158_/A _6253_/C _6075_/C _6075_/D vssd2 vssd2 vccd2 vccd2 _5884_/X sky130_fd_sc_hd__and4_1
X_4835_ _4762_/A _4761_/B _4759_/Y vssd2 vssd2 vccd2 vccd2 _4837_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_269 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7623_ _7627_/A vssd2 vssd2 vccd2 vccd2 _7623_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4044__B _4044_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4766_ _4841_/A _4766_/B vssd2 vssd2 vccd2 vccd2 _4767_/B sky130_fd_sc_hd__or2_2
XFILLER_0_7_355 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__7636__A _7641_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7554_ _7563_/A vssd2 vssd2 vccd2 vccd2 _7554_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_483 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6505_ _6505_/A _6505_/B vssd2 vssd2 vccd2 vccd2 _6507_/A sky130_fd_sc_hd__and2_1
X_4697_ _4641_/A _4641_/B _4642_/X vssd2 vssd2 vccd2 vccd2 _4699_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_250 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7485_ _7725_/Q _7453_/Y _7485_/B1 hold319/X vssd2 vssd2 vccd2 vccd2 _7485_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_101_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6436_ _6436_/A _6437_/A _7222_/B vssd2 vssd2 vccd2 vccd2 _6436_/X sky130_fd_sc_hd__and3_1
XANTENNA__4060__A _7764_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_113_385 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_101_547 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6367_ _6368_/A _6368_/B vssd2 vssd2 vccd2 vccd2 _6367_/X sky130_fd_sc_hd__and2_1
XANTENNA__4343__B1 _5042_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5318_ _5318_/A _5318_/B vssd2 vssd2 vccd2 vccd2 _5320_/B sky130_fd_sc_hd__xnor2_1
X_6298_ _6298_/A _6298_/B vssd2 vssd2 vccd2 vccd2 _6299_/B sky130_fd_sc_hd__xnor2_2
Xhold13 hold13/A vssd2 vssd2 vccd2 vccd2 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7826_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5249_ _5250_/B _5194_/Y _5249_/C _5249_/D vssd2 vssd2 vccd2 vccd2 _5249_/X sky130_fd_sc_hd__and4bb_1
Xhold24 hold24/A vssd2 vssd2 vccd2 vccd2 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd2 vssd2 vccd2 vccd2 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd2 vssd2 vccd2 vccd2 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd2 vssd2 vccd2 vccd2 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd2 vssd2 vccd2 vccd2 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd2 vssd2 vccd2 vccd2 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_648 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_97_125 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_97_169 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_78_350 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_66_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_109_625 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_66_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_109_669 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_81_526 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7546__A _7563_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_19_472 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_46_291 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_261 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_34_464 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_104_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_61_294 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6874__A2 _7294_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_21_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_309 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_57_534 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_29_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XTAP_1092 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_375 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_72_537 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_72_515 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_44_206 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4620_ _4619_/A _4619_/B _4619_/C vssd2 vssd2 vccd2 vccd2 _4621_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_113_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_52_261 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_4_358 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_13_615 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
X_4551_ _4551_/A _4551_/B _4551_/C vssd2 vssd2 vccd2 vccd2 _4552_/B sky130_fd_sc_hd__nand3_1
X_7270_ _7270_/A _7270_/B vssd2 vssd2 vccd2 vccd2 _7271_/B sky130_fd_sc_hd__and2_1
Xhold516 la_data_in[32] vssd2 vssd2 vccd2 vccd2 hold37/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold505 hold11/X vssd2 vssd2 vccd2 vccd2 input3/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_648 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4482_ _4482_/A _4482_/B vssd2 vssd2 vccd2 vccd2 _4484_/A sky130_fd_sc_hd__and2_1
Xhold527 hold60/X vssd2 vssd2 vccd2 vccd2 _7862_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 input25/X vssd2 vssd2 vccd2 vccd2 hold56/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 hold71/X vssd2 vssd2 vccd2 vccd2 input15/A sky130_fd_sc_hd__dlygate4sd3_1
X_6221_ _6158_/A _6510_/B _5751_/Y _7850_/Q vssd2 vssd2 vccd2 vccd2 _6221_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_110_333 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_810 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _6510_/A _6152_/B _6152_/C _6281_/C vssd2 vssd2 vccd2 vccd2 _6152_/X sky130_fd_sc_hd__and4_2
XFILLER_0_40_489 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_110_377 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5103_ _5104_/A _5104_/B vssd2 vssd2 vccd2 vccd2 _5178_/A sky130_fd_sc_hd__nor2_1
XTAP_843 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6082_/A _6571_/A _6082_/C vssd2 vssd2 vccd2 vccd2 _6084_/B sky130_fd_sc_hd__a21o_1
XTAP_876 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5142__C _5142_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5034_ _5160_/A _5033_/C _5033_/A vssd2 vssd2 vccd2 vccd2 _5035_/C sky130_fd_sc_hd__o21ai_1
XTAP_898 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_103 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_18_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_79_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6985_ _7047_/A _7222_/C vssd2 vssd2 vccd2 vccd2 _6988_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4055__A _4898_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5936_ _6510_/A _5936_/B _5936_/C vssd2 vssd2 vccd2 vccd2 _5947_/A sky130_fd_sc_hd__and3_1
XFILLER_0_48_567 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_90_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5867_ _7807_/D _5868_/B _5866_/Y vssd2 vssd2 vccd2 vccd2 _5867_/X sky130_fd_sc_hd__o21ba_1
X_7606_ _7627_/A vssd2 vssd2 vccd2 vccd2 _7606_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7366__A _7436_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_105_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6553__A1 _5991_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4818_ _4818_/A _4818_/B vssd2 vssd2 vccd2 vccd2 _4819_/B sky130_fd_sc_hd__xnor2_4
X_5798_ _5798_/A _5798_/B _5798_/C _5798_/D vssd2 vssd2 vccd2 vccd2 _5798_/Y sky130_fd_sc_hd__nor4_1
XFILLER_0_105_149 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_90_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4749_ _4749_/A _4749_/B vssd2 vssd2 vccd2 vccd2 _4752_/A sky130_fd_sc_hd__xnor2_1
X_7537_ _7561_/A vssd2 vssd2 vccd2 vccd2 _7537_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_453 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_71_592 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_43_294 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7468_ _7708_/Q _7483_/A2 _7483_/B1 hold323/X vssd2 vssd2 vccd2 vccd2 _7468_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_31_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6419_ _6419_/A _6419_/B vssd2 vssd2 vccd2 vccd2 _6421_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_478 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_113_193 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_101_355 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7399_ _7440_/A _7399_/B vssd2 vssd2 vccd2 vccd2 _7668_/D sky130_fd_sc_hd__and2_1
XFILLER_0_101_377 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_98_412 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_98_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_58_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_85_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_534 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_142 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_131 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_120 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_93_161 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XPHY_175 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_164 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_153 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_54_537 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_186 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6544__A1 _5778_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_54_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_26_239 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_22_401 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_34_250 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_78_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_22_434 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_33 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_89_401 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_89_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6355__A _6668_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6770_ _7034_/A _7033_/A vssd2 vssd2 vccd2 vccd2 _6771_/B sky130_fd_sc_hd__nor2_1
XPHY_0 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3982_ _4068_/B _3982_/B _4022_/B _4162_/B vssd2 vssd2 vccd2 vccd2 _4070_/D sky130_fd_sc_hd__nor4_2
XFILLER_0_9_439 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5721_ _5992_/B _5781_/B vssd2 vssd2 vccd2 vccd2 _5845_/B sky130_fd_sc_hd__or2_1
XFILLER_0_57_397 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6802__B _6973_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_84_194 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_72_356 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5652_ _7313_/A _6474_/A vssd2 vssd2 vccd2 vccd2 _6396_/B sky130_fd_sc_hd__nor2_1
X_4603_ _4603_/A _4603_/B vssd2 vssd2 vccd2 vccd2 _4605_/B sky130_fd_sc_hd__xor2_2
X_5583_ _5583_/A _5583_/B vssd2 vssd2 vccd2 vccd2 _6629_/B sky130_fd_sc_hd__and2_1
Xhold302 hold302/A vssd2 vssd2 vccd2 vccd2 la_data_out[22] sky130_fd_sc_hd__buf_12
X_7322_ _7308_/B _7307_/Y _7321_/X vssd2 vssd2 vccd2 vccd2 _7324_/B sky130_fd_sc_hd__o21ai_4
X_4534_ _4534_/A _4534_/B vssd2 vssd2 vccd2 vccd2 _4535_/B sky130_fd_sc_hd__xor2_2
Xhold313 hold666/X vssd2 vssd2 vccd2 vccd2 hold667/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 _7744_/Q vssd2 vssd2 vccd2 vccd2 hold335/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 _7468_/X vssd2 vssd2 vccd2 vccd2 _7708_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_456 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_40_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_111_653 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_110_141 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4465_ _4465_/A _4465_/B vssd2 vssd2 vccd2 vccd2 _4467_/B sky130_fd_sc_hd__xnor2_1
X_7253_ _7253_/A _7253_/B _7253_/C _7253_/D vssd2 vssd2 vccd2 vccd2 _7254_/B sky130_fd_sc_hd__or4_1
Xhold346 _7481_/X vssd2 vssd2 vccd2 vccd2 _7721_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 hold681/X vssd2 vssd2 vccd2 vccd2 _7771_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 _7687_/Q vssd2 vssd2 vccd2 vccd2 hold357/X sky130_fd_sc_hd__dlygate4sd3_1
X_6204_ _6707_/A _6973_/B vssd2 vssd2 vccd2 vccd2 _6206_/A sky130_fd_sc_hd__or2_1
X_7184_ _7144_/A _7146_/B _7144_/B vssd2 vssd2 vccd2 vccd2 _7186_/B sky130_fd_sc_hd__o21ba_1
X_4396_ _4338_/A _4337_/A _4337_/B vssd2 vssd2 vccd2 vccd2 _4404_/A sky130_fd_sc_hd__a21boi_4
Xhold379 _7649_/Q vssd2 vssd2 vccd2 vccd2 hold379/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_297 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6135_ _6572_/B vssd2 vssd2 vccd2 vccd2 _6657_/B sky130_fd_sc_hd__inv_2
XTAP_651 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _6068_/A _6068_/B _7336_/A vssd2 vssd2 vccd2 vccd2 _6067_/B sky130_fd_sc_hd__o21a_1
XTAP_662 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5017_ _5017_/A _5017_/B vssd2 vssd2 vccd2 vccd2 _5021_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__6265__A _6634_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_95_404 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_67_117 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6968_ _6908_/A _6908_/B _6903_/X vssd2 vssd2 vccd2 vccd2 _6969_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_331 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6899_ _6900_/A _6900_/B vssd2 vssd2 vccd2 vccd2 _6899_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_526 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_36_537 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5919_ _6157_/A _6253_/B _6191_/C _6191_/D vssd2 vssd2 vccd2 vccd2 _5923_/A sky130_fd_sc_hd__and4_1
XFILLER_0_75_194 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_91_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_90_153 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5328__B _5528_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_90_197 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4001__A2 _4809_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_7_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__3799__A _7767_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_98_253 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6214__B1 _6150_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_58_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_104_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_39_353 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4776__B1 _5076_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_13_35 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_526 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_82_654 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_81_120 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__6517__A1 _6668_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_6_409 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_89_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_81_164 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_42_507 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_22_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_1_158 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4250_ _7771_/Q _4160_/B _4057_/X _4268_/A _4249_/X vssd2 vssd2 vccd2 vccd2 _4250_/X
+ sky130_fd_sc_hd__a221o_1
X_4181_ _4181_/A _4181_/B vssd2 vssd2 vccd2 vccd2 _4183_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_54 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5404__D _5498_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7871_ _7878_/CLK _7871_/D _7630_/Y vssd2 vssd2 vccd2 vccd2 _7871_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5008__B2 _5168_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5008__A1 _5207_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6822_ _6822_/A _6822_/B vssd2 vssd2 vccd2 vccd2 _6825_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_85_470 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6753_ _6753_/A _6753_/B vssd2 vssd2 vccd2 vccd2 _6754_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_64_109 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_57_172 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_9_236 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3965_ _3965_/A _4033_/C vssd2 vssd2 vccd2 vccd2 _3965_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85_492 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6684_ _6684_/A _6684_/B vssd2 vssd2 vccd2 vccd2 _6685_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__4333__A _4810_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5704_ _7885_/Q _5704_/B vssd2 vssd2 vccd2 vccd2 _6588_/B sky130_fd_sc_hd__xor2_4
X_3896_ _4814_/A _4458_/C _4141_/C _3896_/D vssd2 vssd2 vccd2 vccd2 _3904_/B sky130_fd_sc_hd__or4_2
XFILLER_0_73_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_73_665 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_72_153 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5635_ _5645_/B _7859_/Q _7860_/Q _5641_/B vssd2 vssd2 vccd2 vccd2 _5638_/C sky130_fd_sc_hd__a211o_1
XFILLER_0_85_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_45_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_79_61 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold110 wbs_adr_i[2] vssd2 vssd2 vccd2 vccd2 input72/A sky130_fd_sc_hd__dlygate4sd3_1
X_5566_ _5566_/A _5566_/B vssd2 vssd2 vccd2 vccd2 _7755_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__3891__B _7763_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7305_ _7303_/A _7303_/B _7303_/C vssd2 vssd2 vccd2 vccd2 _7306_/B sky130_fd_sc_hd__o21a_1
X_4517_ _4517_/A _4517_/B vssd2 vssd2 vccd2 vccd2 _4535_/A sky130_fd_sc_hd__xor2_2
Xhold143 hold385/X vssd2 vssd2 vccd2 vccd2 _7766_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 input97/X vssd2 vssd2 vccd2 vccd2 hold121/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 wbs_adr_i[26] vssd2 vssd2 vccd2 vccd2 input68/A sky130_fd_sc_hd__dlygate4sd3_1
X_5497_ _5550_/A _5528_/A _5498_/D _5498_/A vssd2 vssd2 vccd2 vccd2 _5499_/A sky130_fd_sc_hd__o22ai_1
X_7236_ _7236_/A _7236_/B vssd2 vssd2 vccd2 vccd2 _7239_/B sky130_fd_sc_hd__xor2_1
X_4448_ _4448_/A _4448_/B vssd2 vssd2 vccd2 vccd2 _4449_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__7484__A2 _7454_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold154 _7353_/X vssd2 vssd2 vccd2 vccd2 _7354_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_670 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold165 _7421_/X vssd2 vssd2 vccd2 vccd2 _7422_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _7423_/X vssd2 vssd2 vccd2 vccd2 _7424_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 input91/X vssd2 vssd2 vccd2 vccd2 hold187/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold198 hold396/X vssd2 vssd2 vccd2 vccd2 _7772_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7167_ _7167_/A _7167_/B vssd2 vssd2 vccd2 vccd2 _7168_/B sky130_fd_sc_hd__nor2_1
X_4379_ _4708_/A _5220_/A vssd2 vssd2 vccd2 vccd2 _4393_/A sky130_fd_sc_hd__nor2_1
X_6118_ _6115_/Y _6116_/X _6055_/B _6057_/B vssd2 vssd2 vccd2 vccd2 _6119_/C sky130_fd_sc_hd__o211a_1
XANTENNA__6707__B _7255_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7098_ _7098_/A _7098_/B vssd2 vssd2 vccd2 vccd2 _7100_/A sky130_fd_sc_hd__nand2_1
XTAP_470 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _6049_/A _6049_/B _6049_/C vssd2 vssd2 vccd2 vccd2 _6051_/B sky130_fd_sc_hd__nand3_1
XTAP_1614 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_68_415 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XTAP_1625 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_610 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_49_673 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_36_312 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_76_481 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_63_131 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_36_356 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_233 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__7554__A _7563_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_24_529 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_106_277 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_51_348 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_461 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7475__A2 _7483_/A2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_102_483 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_99_540 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_99_573 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_86_289 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_74_418 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_55_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7163__A1 _7045_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_54_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__3992__A _4598_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_42_348 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5420_ _5421_/A _5420_/B _5421_/B vssd2 vssd2 vccd2 vccd2 _5422_/B sky130_fd_sc_hd__and3_1
X_5351_ _5301_/A _5301_/B _5299_/X vssd2 vssd2 vccd2 vccd2 _5353_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__4600__B _5374_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_49_53 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5282_ _5404_/A _5406_/A _5498_/A _5431_/A vssd2 vssd2 vccd2 vccd2 _5284_/A sky130_fd_sc_hd__o22a_1
XFILLER_0_10_234 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7466__A2 _7454_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4302_ _4360_/A _4302_/B vssd2 vssd2 vccd2 vccd2 _4304_/B sky130_fd_sc_hd__nand2_1
X_7021_ _6847_/A _6847_/B _6964_/B _6963_/B _6963_/A vssd2 vssd2 vccd2 vccd2 _7024_/B
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_10_267 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5477__A1 _4893_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4233_ _4234_/A _4234_/B vssd2 vssd2 vccd2 vccd2 _4293_/A sky130_fd_sc_hd__nand2b_1
X_4164_ _4814_/A _4214_/C _4164_/C vssd2 vssd2 vccd2 vccd2 _4164_/X sky130_fd_sc_hd__or3_1
XANTENNA__4328__A _4328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4095_ _4095_/A _4096_/B vssd2 vssd2 vccd2 vccd2 _7729_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__5431__B _5431_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_77_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_77_212 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7639__A _7641_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_81_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7854_ _7854_/CLK _7854_/D _7613_/Y vssd2 vssd2 vccd2 vccd2 _7854_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_278 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_65_429 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7785_ _7787_/CLK _7785_/D _7544_/Y vssd2 vssd2 vccd2 vccd2 _7785_/Q sky130_fd_sc_hd__dfrtp_4
X_6805_ _6804_/A _6876_/A _6804_/C vssd2 vssd2 vccd2 vccd2 _6806_/C sky130_fd_sc_hd__a21o_1
X_6736_ _5890_/A _5890_/B _6664_/A _7222_/B _7294_/C vssd2 vssd2 vccd2 vccd2 _6737_/B
+ sky130_fd_sc_hd__o2111a_1
X_4997_ _4997_/A _4997_/B vssd2 vssd2 vccd2 vccd2 _5133_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_61_613 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3948_ _3941_/X _3947_/X _4315_/C vssd2 vssd2 vccd2 vccd2 _3948_/X sky130_fd_sc_hd__o21a_1
X_6667_ _6667_/A _6667_/B vssd2 vssd2 vccd2 vccd2 _6677_/A sky130_fd_sc_hd__xnor2_2
X_3879_ _3879_/A vssd2 vssd2 vccd2 vccd2 _3880_/D sky130_fd_sc_hd__inv_2
XANTENNA__4998__A _5548_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7374__A _7452_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_33_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6598_ _6599_/A _6599_/B vssd2 vssd2 vccd2 vccd2 _6598_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_14_551 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5618_ _7844_/Q _6191_/D vssd2 vssd2 vccd2 vccd2 _5618_/X sky130_fd_sc_hd__and2_1
XFILLER_0_103_225 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4510__B _5099_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5549_ _5549_/A _5549_/B vssd2 vssd2 vccd2 vccd2 _7754_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__7457__A2 _7454_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7219_ _7336_/A _7219_/B vssd2 vssd2 vccd2 vccd2 _7220_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_96_521 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_68_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4443__A2 _4965_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1433 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_289 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1499 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_248 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_36_120 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_64_451 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_37_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_107_553 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_91_281 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_64_495 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_36_175 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_107_586 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_101_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_10_36 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_24_348 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_24_359 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_86_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_32_381 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6628__A _6670_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_554 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_87_543 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4920_ _4920_/A _4920_/B vssd2 vssd2 vccd2 vccd2 _4923_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_88 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6082__B _6571_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4851_ _4845_/A _4845_/B _4842_/A vssd2 vssd2 vccd2 vccd2 _4925_/A sky130_fd_sc_hd__a21boi_4
XANTENNA__7178__B _7255_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_289 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3802_ _6283_/A vssd2 vssd2 vccd2 vccd2 _6358_/A sky130_fd_sc_hd__inv_2
X_7570_ _7613_/A vssd2 vssd2 vccd2 vccd2 _7570_/Y sky130_fd_sc_hd__inv_2
X_4782_ _5210_/A _4782_/B _5099_/A _4965_/B vssd2 vssd2 vccd2 vccd2 _4783_/B sky130_fd_sc_hd__or4_1
X_6521_ _6442_/A _6442_/B _6440_/X vssd2 vssd2 vccd2 vccd2 _6523_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_70_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6452_ _6452_/A _6452_/B vssd2 vssd2 vccd2 vccd2 _6453_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_359 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_42_134 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_30_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5403_ _5498_/A _5468_/A _5498_/D _5404_/A vssd2 vssd2 vccd2 vccd2 _5403_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_42_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_113_567 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6383_ _6384_/B _6384_/A vssd2 vssd2 vccd2 vccd2 _6457_/A sky130_fd_sc_hd__nand2b_1
X_5334_ _5379_/A _5334_/B vssd2 vssd2 vccd2 vccd2 _5335_/B sky130_fd_sc_hd__nand2_1
X_5265_ _5266_/A _5266_/B vssd2 vssd2 vccd2 vccd2 _5265_/Y sky130_fd_sc_hd__nand2_1
X_5196_ _5250_/B _5130_/B _5125_/X vssd2 vssd2 vccd2 vccd2 _5197_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_48_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4216_ _4315_/C _3943_/X _4215_/X _4160_/B _4162_/A vssd2 vssd2 vccd2 vccd2 _4216_/X
+ sky130_fd_sc_hd__a32o_1
X_7004_ _7004_/A _7004_/B vssd2 vssd2 vccd2 vccd2 _7005_/B sky130_fd_sc_hd__xor2_1
XANTENNA__6257__B _7051_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5870__A1 _7336_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4147_ _7764_/Q _4809_/B vssd2 vssd2 vccd2 vccd2 _4147_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_78_521 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4078_ _7762_/Q _4809_/B _3892_/B _4076_/X _4073_/X vssd2 vssd2 vccd2 vccd2 _4078_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_92_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6273__A _6581_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_78_554 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7837_ _7838_/CLK _7837_/D _7596_/Y vssd2 vssd2 vccd2 vccd2 _7837_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_557 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_65_248 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7768_ _7768_/CLK _7768_/D _7527_/Y vssd2 vssd2 vccd2 vccd2 _7768_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_73_270 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6719_ _6719_/A _6719_/B vssd2 vssd2 vccd2 vccd2 _6721_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_495 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_46_473 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7699_ _7798_/CLK _7699_/D vssd2 vssd2 vccd2 vccd2 _7699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_454 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_443 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5617__A _7845_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_104_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_61_476 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_21_318 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_104_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6638__B1 _7143_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout250 _4522_/C vssd2 vssd2 vccd2 vccd2 _4454_/B sky130_fd_sc_hd__clkbuf_8
Xfanout261 _7851_/Q vssd2 vssd2 vccd2 vccd2 _6283_/A sky130_fd_sc_hd__buf_4
Xfanout283 _7563_/A vssd2 vssd2 vccd2 vccd2 _7561_/A sky130_fd_sc_hd__buf_8
Xfanout272 _7772_/Q vssd2 vssd2 vccd2 vccd2 _4268_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6810__B1 _7294_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_84_513 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1241 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_418 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1263 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_557 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1252 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1296 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_21_35 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_114_309 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_107_361 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4431__A _4598_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_21_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_21_79 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_24_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_97_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_20_351 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5050_ _5051_/A _5051_/B vssd2 vssd2 vccd2 vccd2 _5050_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4444__C_N _5030_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4104__A1 _4268_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4001_ _7761_/Q _4809_/B _4146_/B _7762_/Q vssd2 vssd2 vccd2 vccd2 _4001_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_46_76 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5952_ _5952_/A _5952_/B _5952_/C vssd2 vssd2 vccd2 vccd2 _5956_/A sky130_fd_sc_hd__and3_1
XANTENNA__6801__B1 _7099_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6093__A _6093_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_75_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5080__A2 _5406_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4903_ _4903_/A _4903_/B vssd2 vssd2 vccd2 vccd2 _4904_/B sky130_fd_sc_hd__xor2_4
X_5883_ _5883_/A _5883_/B _5883_/C _5883_/D vssd2 vssd2 vccd2 vccd2 _6424_/B sky130_fd_sc_hd__or4_4
XFILLER_0_90_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4834_ _4834_/A _4834_/B vssd2 vssd2 vccd2 vccd2 _4837_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_568 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7622_ _7627_/A vssd2 vssd2 vccd2 vccd2 _7622_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_90_538 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4765_ _4765_/A _4765_/B vssd2 vssd2 vccd2 vccd2 _4766_/B sky130_fd_sc_hd__and2_1
XFILLER_0_7_345 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7553_ _7557_/A vssd2 vssd2 vccd2 vccd2 _7553_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_473 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6504_ _6812_/A _6812_/B _7140_/A _7237_/A vssd2 vssd2 vccd2 vccd2 _6505_/B sky130_fd_sc_hd__or4_1
XFILLER_0_43_454 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_16_668 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA_fanout219_A _4628_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4696_ _4687_/Y _4691_/B _4686_/A vssd2 vssd2 vccd2 vccd2 _4768_/A sky130_fd_sc_hd__o21ai_2
X_7484_ _7724_/Q _7454_/C _7485_/B1 hold321/X vssd2 vssd2 vccd2 vccd2 _7484_/X sky130_fd_sc_hd__a22o_1
X_6435_ _6436_/A _7222_/B vssd2 vssd2 vccd2 vccd2 _6437_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_126 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_101_515 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6366_ _6668_/A _7094_/A _6290_/B _6288_/X vssd2 vssd2 vccd2 vccd2 _6368_/B sky130_fd_sc_hd__a31o_1
XANTENNA__4343__A1 _4044_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_101_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6268__A _6707_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5317_ _5431_/A _5550_/A vssd2 vssd2 vccd2 vccd2 _5318_/B sky130_fd_sc_hd__nor2_1
X_6297_ _6298_/B _6298_/A vssd2 vssd2 vccd2 vccd2 _6297_/Y sky130_fd_sc_hd__nand2b_1
Xhold14 hold14/A vssd2 vssd2 vccd2 vccd2 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd2 vssd2 vccd2 vccd2 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
X_5248_ _5248_/A _5248_/B vssd2 vssd2 vccd2 vccd2 _5447_/A sky130_fd_sc_hd__xor2_1
Xhold36 hold36/A vssd2 vssd2 vccd2 vccd2 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd2 vssd2 vccd2 vccd2 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd2 vssd2 vccd2 vccd2 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
X_5179_ _4172_/Y _5550_/B _5233_/A _5178_/Y vssd2 vssd2 vccd2 vccd2 _5182_/A sky130_fd_sc_hd__o22a_1
Xhold58 hold58/A vssd2 vssd2 vccd2 vccd2 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_137 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7099__A _7145_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_78_362 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_93_376 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6020__A1 _7850_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_19_495 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_34_421 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4251__A _4656_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_22_627 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_34_487 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5531__B1 _5550_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_100_570 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_107_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_89_649 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_16_24 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_97_671 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_57_513 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__3968__C _7766_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1082 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_387 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1093 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3984__B _5030_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_65_590 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5257__A _5257_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_37_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_106_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_80_571 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_25_465 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4550_ _4551_/B _4551_/C _4551_/A vssd2 vssd2 vccd2 vccd2 _4619_/B sky130_fd_sc_hd__a21o_1
Xhold517 hold37/X vssd2 vssd2 vccd2 vccd2 input26/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold506 input3/X vssd2 vssd2 vccd2 vccd2 hold12/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_498 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4481_ _4480_/A _4480_/B _4480_/C vssd2 vssd2 vccd2 vccd2 _4482_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_110_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6220_ _6093_/A _6281_/B _6152_/C _6253_/A vssd2 vssd2 vccd2 vccd2 _6220_/X sky130_fd_sc_hd__a22o_1
Xhold528 la_data_in[24] vssd2 vssd2 vccd2 vccd2 hold53/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 hold56/X vssd2 vssd2 vccd2 vccd2 _7870_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap247 _4006_/B vssd2 vssd2 vccd2 vccd2 _4893_/B sky130_fd_sc_hd__buf_4
XANTENNA__4325__B2 _7768_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4325__A1 _4162_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_110_345 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6151_ _5816_/A _5816_/B _6571_/C vssd2 vssd2 vccd2 vccd2 _6164_/A sky130_fd_sc_hd__a21boi_2
XTAP_800 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_389 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5102_ _5220_/A _5222_/A _5041_/X _5043_/B vssd2 vssd2 vccd2 vccd2 _5104_/B sky130_fd_sc_hd__o31a_1
XTAP_844 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6082_/A _6571_/A _6082_/C vssd2 vssd2 vccd2 vccd2 _6144_/A sky130_fd_sc_hd__and3_1
XTAP_877 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5142__D _5498_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5033_ _5033_/A _5160_/A _5033_/C vssd2 vssd2 vccd2 vccd2 _5035_/B sky130_fd_sc_hd__or3_1
XTAP_899 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_74 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4336__A _4863_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_fanout169_A _6705_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5589__B1 _5645_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6984_ _6928_/A _6928_/B _6926_/Y vssd2 vssd2 vccd2 vccd2 _7003_/A sky130_fd_sc_hd__a21oi_1
X_5935_ _6100_/D _6587_/B _5938_/C _5935_/D vssd2 vssd2 vccd2 vccd2 _5935_/X sky130_fd_sc_hd__and4_1
XANTENNA__4055__B _4882_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5866_ _5917_/A _5866_/B vssd2 vssd2 vccd2 vccd2 _5866_/Y sky130_fd_sc_hd__nand2_1
X_4817_ _4818_/A _4818_/B vssd2 vssd2 vccd2 vccd2 _4817_/X sky130_fd_sc_hd__and2b_1
X_7605_ _7627_/A vssd2 vssd2 vccd2 vccd2 _7605_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_643 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_8_632 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6553__A2 _5993_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_8_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_7_153 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_28_270 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5797_ _7841_/Q _7313_/A _6398_/B _7842_/Q vssd2 vssd2 vccd2 vccd2 _5798_/D sky130_fd_sc_hd__a22o_1
X_4748_ _4748_/A _4748_/B vssd2 vssd2 vccd2 vccd2 _4749_/B sky130_fd_sc_hd__xnor2_1
X_7536_ _7557_/A vssd2 vssd2 vccd2 vccd2 _7536_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_465 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_114_651 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4679_ _4679_/A _4679_/B vssd2 vssd2 vccd2 vccd2 _4681_/B sky130_fd_sc_hd__xnor2_1
X_7467_ _7707_/Q _7454_/C _7485_/B1 hold233/X vssd2 vssd2 vccd2 vccd2 _7467_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_113_161 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6418_ _6855_/A _7037_/A vssd2 vssd2 vccd2 vccd2 _6419_/B sky130_fd_sc_hd__nor2_1
XANTENNA__7382__A _7452_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4316__A1 _7768_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4316__B2 _4162_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_101_345 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7398_ hold172/X _7668_/Q _7418_/S vssd2 vssd2 vccd2 vccd2 _7398_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_101_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6349_ _6581_/A _6989_/A vssd2 vssd2 vccd2 vccd2 _6354_/A sky130_fd_sc_hd__nor2_1
XANTENNA__5006__A2_N _5431_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_79_671 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_78_181 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_39_524 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_94_641 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XPHY_143 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_132 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_121 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_110 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7557__A _7557_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_39_557 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_176 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_165 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_154 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_66_398 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_66_365 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_54_516 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_198 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_187 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_81_346 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_81_324 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6544__A2 _5786_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_19_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_22_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_94_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6355__B _7197_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_77_608 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4156__A _4747_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_57_310 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_43_44 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XPHY_1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3981_ _3930_/X _3980_/X _3979_/X _3969_/X _3948_/X vssd2 vssd2 vccd2 vccd2 _3981_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_43_99 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5720_ _7876_/Q _5720_/B vssd2 vssd2 vccd2 vccd2 _5781_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_72_313 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_72_302 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_45_527 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_45_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6802__C _7237_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_17_229 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5651_ _5811_/B _5811_/C vssd2 vssd2 vccd2 vccd2 _5835_/D sky130_fd_sc_hd__nor2_1
X_4602_ _4603_/A _4603_/B vssd2 vssd2 vccd2 vccd2 _4672_/A sky130_fd_sc_hd__nand2_1
X_5582_ _7867_/Q _7868_/Q vssd2 vssd2 vccd2 vccd2 _5583_/B sky130_fd_sc_hd__nor2_2
X_7321_ _7308_/A _7306_/A _7306_/B vssd2 vssd2 vccd2 vccd2 _7321_/X sky130_fd_sc_hd__o21ba_1
X_4533_ _4534_/A _4534_/B vssd2 vssd2 vccd2 vccd2 _4533_/X sky130_fd_sc_hd__and2_1
XFILLER_0_13_435 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold303 hold656/X vssd2 vssd2 vccd2 vccd2 hold657/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_109 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold314 hold314/A vssd2 vssd2 vccd2 vccd2 la_data_out[11] sky130_fd_sc_hd__buf_12
X_7252_ _7253_/B _7253_/C _7253_/D _7253_/A vssd2 vssd2 vccd2 vccd2 _7252_/X sky130_fd_sc_hd__o22a_1
XANTENNA__7406__S _7418_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold325 _7741_/Q vssd2 vssd2 vccd2 vccd2 hold325/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6203_ _6636_/A _7037_/A vssd2 vssd2 vccd2 vccd2 _6208_/A sky130_fd_sc_hd__nor2_1
X_4464_ _4462_/X _4464_/B vssd2 vssd2 vccd2 vccd2 _4465_/B sky130_fd_sc_hd__nand2b_1
Xhold369 _7669_/Q vssd2 vssd2 vccd2 vccd2 hold369/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 _7747_/Q vssd2 vssd2 vccd2 vccd2 hold347/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _7472_/X vssd2 vssd2 vccd2 vccd2 _7712_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 _7663_/Q vssd2 vssd2 vccd2 vccd2 hold358/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_276 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_111_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_110_153 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_68_96 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7183_ _7259_/A _7183_/B vssd2 vssd2 vccd2 vccd2 _7186_/A sky130_fd_sc_hd__and2_1
X_4395_ _4344_/A _4344_/B _4345_/B _4345_/A vssd2 vssd2 vccd2 vccd2 _4405_/A sky130_fd_sc_hd__a22o_2
XFILLER_0_110_197 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_630 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _6130_/X _6131_/X _6133_/X _6075_/C vssd2 vssd2 vccd2 vccd2 _6572_/B sky130_fd_sc_hd__o31ai_4
XANTENNA__6546__A _6707_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6065_ _6065_/A _6065_/B vssd2 vssd2 vccd2 vccd2 _6067_/A sky130_fd_sc_hd__xnor2_1
XTAP_663 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _5328_/A _5366_/A vssd2 vssd2 vccd2 vccd2 _5017_/B sky130_fd_sc_hd__nor2_1
XANTENNA_fanout286_A _7629_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_30_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XTAP_696 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6265__B _6571_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4066__A _4268_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6967_ _6967_/A _6967_/B vssd2 vssd2 vccd2 vccd2 _7025_/D sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5918_ _5918_/A _5918_/B vssd2 vssd2 vccd2 vccd2 _7810_/D sky130_fd_sc_hd__xnor2_1
X_6898_ _6830_/A _6830_/B _6828_/Y vssd2 vssd2 vccd2 vccd2 _6900_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_48_376 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_48_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_36_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_90_121 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_8_473 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_8_451 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5849_ _7842_/Q _6510_/B _6357_/B _7844_/Q vssd2 vssd2 vccd2 vccd2 _5849_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_90_165 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_51_508 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_44_560 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_16_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7519_ _7557_/A vssd2 vssd2 vccd2 vccd2 _7519_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_31_232 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_31_276 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_98_221 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_98_265 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6214__A1 _6664_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6214__B2 _5931_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_438 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_86_427 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_104_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4776__A1 _5011_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4225__B1 _4896_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4776__B2 _4863_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4704__A _4779_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6517__A2 _6430_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_54_324 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_81_143 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7478__B1 _7483_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_22_265 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4180_ _4180_/A _4180_/B vssd2 vssd2 vccd2 vccd2 _4181_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_77_405 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7870_ _7870_/CLK _7870_/D _7629_/Y vssd2 vssd2 vccd2 vccd2 _7870_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5008__A2 _5142_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_77_416 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6821_ _6820_/A _6820_/B _6820_/C vssd2 vssd2 vccd2 vccd2 _6822_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7197__A _7197_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6813__B _7291_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6752_ _6753_/A _6753_/B vssd2 vssd2 vccd2 vccd2 _6752_/Y sky130_fd_sc_hd__nor2_1
X_3964_ _7776_/Q _3964_/B vssd2 vssd2 vccd2 vccd2 _4033_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_18_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_18_527 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6683_ _6684_/A _6684_/B vssd2 vssd2 vccd2 vccd2 _6683_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_72_121 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__4333__B _5099_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_45_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5703_ _7885_/Q _5704_/B vssd2 vssd2 vccd2 vccd2 _6358_/B sky130_fd_sc_hd__xnor2_2
X_3895_ _4267_/D _3996_/B _3895_/C _3895_/D vssd2 vssd2 vccd2 vccd2 _3896_/D sky130_fd_sc_hd__or4_1
XANTENNA__3875__D _4267_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5634_ _7859_/Q _5581_/A _7860_/Q _5645_/B vssd2 vssd2 vccd2 vccd2 _5638_/B sky130_fd_sc_hd__o211ai_2
XFILLER_0_26_560 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7304_ _7304_/A vssd2 vssd2 vccd2 vccd2 _7306_/A sky130_fd_sc_hd__inv_2
Xhold100 _7348_/X vssd2 vssd2 vccd2 vccd2 _7646_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7469__B1 _7483_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5565_ _5549_/A _5548_/B _5548_/A vssd2 vssd2 vccd2 vccd2 _5566_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_73 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4516_ _4516_/A _4516_/B vssd2 vssd2 vccd2 vccd2 _4517_/B sky130_fd_sc_hd__xor2_2
Xhold122 _7404_/X vssd2 vssd2 vccd2 vccd2 _7405_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 _7367_/X vssd2 vssd2 vccd2 vccd2 _7368_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 input72/X vssd2 vssd2 vccd2 vccd2 _7386_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 input68/X vssd2 vssd2 vccd2 vccd2 _7339_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5496_ _5496_/A _5496_/B vssd2 vssd2 vccd2 vccd2 _5500_/A sky130_fd_sc_hd__or2_1
XFILLER_0_41_574 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7235_ _7236_/A _7236_/B vssd2 vssd2 vccd2 vccd2 _7273_/A sky130_fd_sc_hd__nand2_1
X_4447_ _4448_/A _4448_/B vssd2 vssd2 vccd2 vccd2 _4447_/Y sky130_fd_sc_hd__nand2_1
Xhold166 hold388/X vssd2 vssd2 vccd2 vccd2 _7787_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 hold382/X vssd2 vssd2 vccd2 vccd2 _7776_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 hold370/X vssd2 vssd2 vccd2 vccd2 _7782_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7166_ _7166_/A _7166_/B _7166_/C vssd2 vssd2 vccd2 vccd2 _7167_/B sky130_fd_sc_hd__nor3_1
Xhold188 _7392_/X vssd2 vssd2 vccd2 vccd2 _7393_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _7379_/X vssd2 vssd2 vccd2 vccd2 _7380_/B sky130_fd_sc_hd__dlygate4sd3_1
X_6117_ _6055_/B _6057_/B _6115_/Y _6116_/X vssd2 vssd2 vccd2 vccd2 _6119_/B sky130_fd_sc_hd__a211oi_1
XTAP_460 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4378_ _4375_/X _4377_/X _4162_/B vssd2 vssd2 vccd2 vccd2 _5325_/A sky130_fd_sc_hd__o21ai_2
X_7097_ _7143_/A _7143_/B _7222_/B _7294_/C vssd2 vssd2 vccd2 vccd2 _7098_/B sky130_fd_sc_hd__nand4_1
XTAP_482 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _6049_/A _6049_/B _6049_/C vssd2 vssd2 vccd2 vccd2 _6048_/X sky130_fd_sc_hd__and3_1
XTAP_1615 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_83_408 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_64_600 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_48_162 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_63_110 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_63_143 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_106_289 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_32_541 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_451 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_102_495 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_102_473 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7570__A _7613_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4694__B1 _4693_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4446__B1 _4965_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_99_552 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_59_416 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4434__A _4863_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_24_68 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_27_302 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_39_151 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_82_441 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_40_12 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7163__A2 _7291_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_42_316 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__3992__B _4747_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_27_379 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_23_530 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5350_ _5395_/B _5350_/B vssd2 vssd2 vccd2 vccd2 _5353_/A sky130_fd_sc_hd__and2_2
X_5281_ _5281_/A _5281_/B vssd2 vssd2 vccd2 vccd2 _5289_/A sky130_fd_sc_hd__xnor2_2
X_4301_ _4301_/A _4303_/D vssd2 vssd2 vccd2 vccd2 _4302_/B sky130_fd_sc_hd__nand2_1
XANTENNA__6674__A1 _6668_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7020_ _7081_/B _7020_/B vssd2 vssd2 vccd2 vccd2 _7024_/A sky130_fd_sc_hd__nor2_2
X_4232_ _4232_/A _4232_/B vssd2 vssd2 vccd2 vccd2 _4234_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_65_42 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4163_ _4268_/A _4214_/C vssd2 vssd2 vccd2 vccd2 _4163_/Y sky130_fd_sc_hd__nand2_1
X_4094_ _4094_/A _4189_/B vssd2 vssd2 vccd2 vccd2 _4096_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__5634__C1 _5645_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7853_ _7854_/CLK _7853_/D _7612_/Y vssd2 vssd2 vccd2 vccd2 _7853_/Q sky130_fd_sc_hd__dfrtp_2
X_4996_ _5128_/A _4996_/B vssd2 vssd2 vccd2 vccd2 _5133_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_65_408 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7784_ _7802_/CLK _7784_/D _7543_/Y vssd2 vssd2 vccd2 vccd2 _7784_/Q sky130_fd_sc_hd__dfrtp_4
X_6804_ _6804_/A _6876_/A _6804_/C vssd2 vssd2 vccd2 vccd2 _6876_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_105_81 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_58_482 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6735_ _6424_/A _6424_/B _7294_/C _7222_/B _6664_/A vssd2 vssd2 vccd2 vccd2 _6737_/A
+ sky130_fd_sc_hd__a32oi_2
X_3947_ _4315_/B _4427_/A _3947_/C vssd2 vssd2 vccd2 vccd2 _3947_/X sky130_fd_sc_hd__and3_1
XFILLER_0_73_452 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_73_485 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6666_ _6873_/A _7237_/A vssd2 vssd2 vccd2 vccd2 _6667_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_45_187 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3878_ _4454_/A _3993_/D vssd2 vssd2 vccd2 vccd2 _3879_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_305 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6597_ _6520_/A _6520_/B _6518_/X vssd2 vssd2 vccd2 vccd2 _6599_/B sky130_fd_sc_hd__a21o_1
X_5617_ _7845_/Q _5620_/B _5630_/B vssd2 vssd2 vccd2 vccd2 _5617_/X sky130_fd_sc_hd__and3_1
XFILLER_0_103_237 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5548_ _5548_/A _5548_/B vssd2 vssd2 vccd2 vccd2 _5549_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_14_563 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_41_360 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_41_393 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_111_281 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7218_ _7326_/A _7326_/B _7326_/C vssd2 vssd2 vccd2 vccd2 _7219_/B sky130_fd_sc_hd__nand3_2
X_5479_ _5480_/A _5480_/B _5480_/C vssd2 vssd2 vccd2 vccd2 _5515_/A sky130_fd_sc_hd__o21ai_1
X_7149_ _7149_/A _7149_/B vssd2 vssd2 vccd2 vccd2 _7152_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__4519__A _4656_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_290 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_533 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1401 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1489 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5069__B _5133_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_107_521 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_51_102 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_101_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_91_293 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_51_135 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_87_522 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4223__C_N _5030_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_99_393 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_87_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_59_235 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4850_ _5455_/A _4997_/A vssd2 vssd2 vccd2 vccd2 _4926_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3801_ _6093_/A vssd2 vssd2 vccd2 vccd2 _6154_/A sky130_fd_sc_hd__inv_2
X_6520_ _6520_/A _6520_/B vssd2 vssd2 vccd2 vccd2 _6523_/A sky130_fd_sc_hd__xnor2_2
X_4781_ _5210_/B _5099_/A _4965_/B _5210_/A vssd2 vssd2 vccd2 vccd2 _4781_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_55_441 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_51_88 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_7_527 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_70_400 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_165 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6451_ _6377_/A _6377_/B _6375_/X vssd2 vssd2 vccd2 vccd2 _6452_/B sky130_fd_sc_hd__a21oi_2
X_6382_ _6307_/A _6307_/B _6305_/Y vssd2 vssd2 vccd2 vccd2 _6384_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_70_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_11_500 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5402_ _5402_/A _5547_/C vssd2 vssd2 vccd2 vccd2 _7750_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_371 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5333_ _5333_/A _5333_/B vssd2 vssd2 vccd2 vccd2 _5379_/B sky130_fd_sc_hd__xor2_2
XANTENNA__7414__S _7418_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_76_52 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5264_ _5315_/B _5374_/B vssd2 vssd2 vccd2 vccd2 _5266_/B sky130_fd_sc_hd__nor2_1
X_5195_ _5195_/A _5195_/B vssd2 vssd2 vccd2 vccd2 _5250_/D sky130_fd_sc_hd__xnor2_4
XFILLER_0_76_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4215_ _4268_/A _4214_/B _4214_/Y vssd2 vssd2 vccd2 vccd2 _4215_/X sky130_fd_sc_hd__a21o_1
X_7003_ _7003_/A _7003_/B vssd2 vssd2 vccd2 vccd2 _7004_/B sky130_fd_sc_hd__xnor2_1
X_4146_ _7765_/Q _4146_/B vssd2 vssd2 vccd2 vccd2 _4146_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_78_511 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6554__A _6556_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4077_ _4326_/B _4268_/D _4074_/X _4200_/B _4328_/A vssd2 vssd2 vccd2 vccd2 _4077_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6273__B _6939_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3897__B _4328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7836_ _7838_/CLK _7836_/D _7595_/Y vssd2 vssd2 vccd2 vccd2 _7836_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_514 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_78_566 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_38_408 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_108_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_93_569 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4979_ _4908_/A _4908_/B _4906_/Y vssd2 vssd2 vccd2 vccd2 _4981_/B sky130_fd_sc_hd__a21o_2
X_7767_ _7802_/CLK _7767_/D _7526_/Y vssd2 vssd2 vccd2 vccd2 _7767_/Q sky130_fd_sc_hd__dfrtp_4
X_6718_ _6718_/A _6718_/B vssd2 vssd2 vccd2 vccd2 _6719_/B sky130_fd_sc_hd__xor2_1
X_7698_ _7798_/CLK _7698_/D vssd2 vssd2 vccd2 vccd2 _7698_/Q sky130_fd_sc_hd__dfxtp_1
X_6649_ _6650_/A _6650_/B vssd2 vssd2 vccd2 vccd2 _6651_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4897__B1 _5528_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_14_360 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6638__A1 _5991_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_41_190 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
Xfanout251 _6069_/A vssd2 vssd2 vccd2 vccd2 _7336_/A sky130_fd_sc_hd__buf_4
Xfanout262 _7851_/Q vssd2 vssd2 vccd2 vccd2 _6074_/A sky130_fd_sc_hd__buf_2
Xfanout273 _7771_/Q vssd2 vssd2 vccd2 vccd2 _4454_/A sky130_fd_sc_hd__buf_4
Xfanout284 _7629_/A vssd2 vssd2 vccd2 vccd2 _7563_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__6464__A _7336_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_511 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__6810__A1 _6424_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6810__B2 _6664_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1231 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_408 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1264 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_71_208 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_107_373 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4431__B _5276_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_24_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_37_496 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_52_477 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_52_455 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_12_319 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_24_179 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_110_516 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_20_385 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4159__A _4454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5262__B _5528_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_46_22 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4000_ _4656_/B _4656_/C vssd2 vssd2 vccd2 vccd2 _4146_/B sky130_fd_sc_hd__nor2_2
X_5951_ _6105_/A _6105_/B _6783_/A _6855_/A vssd2 vssd2 vccd2 vccd2 _5952_/C sky130_fd_sc_hd__or4_1
XANTENNA__6093__B _6152_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6801__B2 _6571_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6801__A1 _6571_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_352 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4902_ _4903_/A _4903_/B vssd2 vssd2 vccd2 vccd2 _4902_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_47_238 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_47_216 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5882_ _7849_/Q _5825_/X _5886_/B _5886_/C _5886_/D vssd2 vssd2 vccd2 vccd2 _5883_/D
+ sky130_fd_sc_hd__a2111o_1
X_4833_ _4833_/A _4833_/B vssd2 vssd2 vccd2 vccd2 _4834_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_249 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7621_ _7627_/A vssd2 vssd2 vccd2 vccd2 _7621_/Y sky130_fd_sc_hd__inv_2
X_4764_ _4765_/A _4765_/B vssd2 vssd2 vccd2 vccd2 _4841_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_7_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7552_ _7557_/A vssd2 vssd2 vccd2 vccd2 _7552_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4040__A1 _7762_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6503_ _6425_/A _7197_/A _6430_/B _5931_/C vssd2 vssd2 vccd2 vccd2 _6505_/A sky130_fd_sc_hd__a22o_1
XANTENNA__4341__B _5030_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7483_ _7723_/Q _7483_/A2 _7483_/B1 hold349/X vssd2 vssd2 vccd2 vccd2 _7483_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4040__B2 _7766_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_43_466 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4695_ _5548_/A _4849_/C vssd2 vssd2 vccd2 vccd2 _4769_/A sky130_fd_sc_hd__or2_1
XFILLER_0_15_157 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6434_ _6253_/A _5713_/Y _5752_/Y _6510_/A _6432_/X vssd2 vssd2 vccd2 vccd2 _7291_/A
+ sky130_fd_sc_hd__o221ai_4
XFILLER_0_30_105 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_101_538 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_87_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6365_ _6365_/A _6365_/B vssd2 vssd2 vccd2 vccd2 _6368_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4343__A2 _4044_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6549__A _6670_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_30_138 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_30_149 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6296_ _6234_/A _6232_/Y _6231_/Y vssd2 vssd2 vccd2 vccd2 _6298_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_11_374 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5316_ _5316_/A _5316_/B vssd2 vssd2 vccd2 vccd2 _5318_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6268__B _7037_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5247_ _5247_/A _5247_/B vssd2 vssd2 vccd2 vccd2 _5254_/A sky130_fd_sc_hd__nor2_2
XANTENNA__7293__A1 _7253_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold26 hold26/A vssd2 vssd2 vccd2 vccd2 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd2 vssd2 vccd2 vccd2 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd2 vssd2 vccd2 vccd2 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ _5178_/A _5178_/B _5178_/C vssd2 vssd2 vccd2 vccd2 _5178_/Y sky130_fd_sc_hd__nor3_1
Xhold59 hold59/A vssd2 vssd2 vccd2 vccd2 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd2 vssd2 vccd2 vccd2 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4129_ _4123_/X _4124_/X _4126_/X _4128_/X _4018_/A vssd2 vssd2 vccd2 vccd2 _4129_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_0_97_149 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7099__B _7099_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_66_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_38_205 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7819_ _7826_/CLK _7819_/D _7578_/Y vssd2 vssd2 vccd2 vccd2 _7819_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_569 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_81_539 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_34_400 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_46_271 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_34_433 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_104_321 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_104_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5531__B2 _5498_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5531__A1 _5550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_107_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7036__A1 _6973_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7036__B2 _6973_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6194__A _6253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_88_127 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_16_36 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_69_374 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4270__A1 _4454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1083 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_569 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1094 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3984__C _4162_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_107_181 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold518 input26/X vssd2 vssd2 vccd2 vccd2 hold38/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold507 hold12/X vssd2 vssd2 vccd2 vccd2 _7882_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap226 _6102_/B vssd2 vssd2 vccd2 vccd2 _6281_/C sky130_fd_sc_hd__buf_6
X_4480_ _4480_/A _4480_/B _4480_/C vssd2 vssd2 vccd2 vccd2 _4482_/A sky130_fd_sc_hd__nand3_1
Xmax_cap215 _6078_/Y vssd2 vssd2 vccd2 vccd2 _6920_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_425 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_40_436 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold529 hold53/X vssd2 vssd2 vccd2 vccd2 input17/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_458 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_110_357 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6150_ _6150_/A _6150_/B vssd2 vssd2 vccd2 vccd2 _6165_/A sky130_fd_sc_hd__nand2_1
XTAP_801 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_43 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5101_ _5101_/A _5101_/B vssd2 vssd2 vccd2 vccd2 _5104_/A sky130_fd_sc_hd__xnor2_1
XTAP_834 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _6550_/A _6973_/B vssd2 vssd2 vccd2 vccd2 _6082_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_57_54 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_867 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _5033_/A _5160_/A _5033_/C vssd2 vssd2 vccd2 vccd2 _5091_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_57_98 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_889 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_20 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7750_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_53 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6983_ _6950_/A _6950_/B _6948_/X vssd2 vssd2 vccd2 vccd2 _7004_/A sky130_fd_sc_hd__a21o_1
X_5934_ _6092_/A _6138_/A vssd2 vssd2 vccd2 vccd2 _5952_/A sky130_fd_sc_hd__nor2_1
X_5865_ _5865_/A _5868_/C vssd2 vssd2 vccd2 vccd2 _5866_/B sky130_fd_sc_hd__or2_1
XFILLER_0_8_611 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_75_377 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7604_ _7627_/A vssd2 vssd2 vccd2 vccd2 _7604_/Y sky130_fd_sc_hd__inv_2
X_4816_ _3904_/A _3904_/B _3904_/C _5528_/B vssd2 vssd2 vccd2 vccd2 _4818_/B sky130_fd_sc_hd__a31oi_4
XFILLER_0_113_81 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5796_ _5586_/B _5584_/Y _5586_/Y _5594_/B _5594_/C vssd2 vssd2 vccd2 vccd2 _6398_/B
+ sky130_fd_sc_hd__o2111a_4
XFILLER_0_16_433 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_71_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_71_550 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4747_ _4747_/A _4748_/A _5528_/A vssd2 vssd2 vccd2 vccd2 _4803_/B sky130_fd_sc_hd__or3_1
X_7535_ _7557_/A vssd2 vssd2 vccd2 vccd2 _7535_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5761__B2 _5736_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_16_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_114_641 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4678_ _4610_/A _4610_/B _4608_/Y vssd2 vssd2 vccd2 vccd2 _4679_/B sky130_fd_sc_hd__a21oi_1
X_7466_ _7706_/Q _7454_/C _7485_/B1 hold245/X vssd2 vssd2 vccd2 vccd2 _7466_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_98_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6417_ _6415_/X _6417_/B vssd2 vssd2 vccd2 vccd2 _6419_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__6279__A _6668_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7397_ _7440_/A _7397_/B vssd2 vssd2 vccd2 vccd2 _7667_/D sky130_fd_sc_hd__and2_1
X_6348_ _6348_/A _6348_/B vssd2 vssd2 vccd2 vccd2 _6373_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_101_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6279_ _6668_/A _7094_/A vssd2 vssd2 vccd2 vccd2 _6290_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5277__B1 _5550_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_98_469 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_66_300 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_100 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_122 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_109_446 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_166 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_155 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_144 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_66_377 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5358__A _5455_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4262__A _7768_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_109_479 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XPHY_199 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_188 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_177 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7573__A _7613_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_81_358 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_62_572 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_22_414 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5504__A1 _5406_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_34_296 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_104_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7257__A1 _7181_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6636__B _7255_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_27_46 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_27_68 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4491__A1 _4893_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4156__B _4896_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_9_408 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XPHY_2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3980_ _7761_/Q _4063_/B _4814_/B vssd2 vssd2 vccd2 vccd2 _3980_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_43_78 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_57_388 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_57_377 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4172__A _5030_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6802__D _7224_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5650_ _6510_/A _5661_/B _5836_/B _5649_/C _5638_/X vssd2 vssd2 vccd2 vccd2 _5650_/X
+ sky130_fd_sc_hd__a41o_1
X_4601_ _4601_/A _4601_/B vssd2 vssd2 vccd2 vccd2 _4603_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_45_539 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_5_625 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5581_ _5581_/A _5581_/B _5581_/C _5581_/D vssd2 vssd2 vccd2 vccd2 _5583_/A sky130_fd_sc_hd__nor4_2
X_4532_ _4532_/A _4532_/B vssd2 vssd2 vccd2 vccd2 _4534_/B sky130_fd_sc_hd__xnor2_2
X_7320_ _7334_/A _7320_/B vssd2 vssd2 vccd2 vccd2 _7324_/A sky130_fd_sc_hd__nand2_2
Xhold304 hold304/A vssd2 vssd2 vccd2 vccd2 la_data_out[29] sky130_fd_sc_hd__buf_12
Xhold315 hold668/X vssd2 vssd2 vccd2 vccd2 hold669/A sky130_fd_sc_hd__dlygate4sd3_1
X_7251_ _7310_/B _7251_/B vssd2 vssd2 vccd2 vccd2 _7832_/D sky130_fd_sc_hd__xnor2_1
X_4463_ _4962_/A _4896_/A _4662_/B _5099_/A vssd2 vssd2 vccd2 vccd2 _4464_/B sky130_fd_sc_hd__or4_1
Xhold326 _7469_/X vssd2 vssd2 vccd2 vccd2 _7709_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_447 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6099__A _6157_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_40_233 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_111_633 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_110_121 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6202_ _6149_/A _6149_/B _6148_/B vssd2 vssd2 vccd2 vccd2 _6210_/A sky130_fd_sc_hd__o21ai_2
Xhold337 _7748_/Q vssd2 vssd2 vccd2 vccd2 hold337/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 _7475_/X vssd2 vssd2 vccd2 vccd2 _7715_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold359 _7648_/Q vssd2 vssd2 vccd2 vccd2 hold359/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_266 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_110_165 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7182_ _7181_/A _7253_/C _7181_/C vssd2 vssd2 vccd2 vccd2 _7183_/B sky130_fd_sc_hd__o21ai_1
X_4394_ _4468_/A _4394_/B vssd2 vssd2 vccd2 vccd2 _4407_/A sky130_fd_sc_hd__and2_2
XTAP_620 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6133_ _6397_/A _5791_/X _5810_/X _6074_/A _6132_/X vssd2 vssd2 vccd2 vccd2 _6133_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_41 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6064_ _6064_/A _6064_/B _6065_/A vssd2 vssd2 vccd2 vccd2 _6311_/A sky130_fd_sc_hd__or3b_1
XTAP_653 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6546__B _7253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5015_ _5013_/X _5015_/B vssd2 vssd2 vccd2 vccd2 _5017_/A sky130_fd_sc_hd__nand2b_1
XTAP_697 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_85 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA_fanout279_A _7450_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA_fanout181_A _6572_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6966_ _6967_/A _6967_/B vssd2 vssd2 vccd2 vccd2 _6966_/X sky130_fd_sc_hd__and2_1
XFILLER_0_95_428 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5917_ _5917_/A _5967_/B vssd2 vssd2 vccd2 vccd2 _5918_/B sky130_fd_sc_hd__xnor2_1
X_6897_ _6897_/A _6897_/B vssd2 vssd2 vccd2 vccd2 _6900_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_63_303 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_48_388 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4082__A _4656_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6281__B _6281_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_91_645 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_8_463 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5848_ _6100_/D _6094_/B _6587_/B vssd2 vssd2 vccd2 vccd2 _6357_/B sky130_fd_sc_hd__and3_2
XFILLER_0_90_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_16_230 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5779_ _7841_/Q _6588_/B _5751_/Y _7842_/Q vssd2 vssd2 vccd2 vccd2 _5779_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_90_177 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4810__A _4810_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_44_572 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7518_ _7524_/A vssd2 vssd2 vccd2 vccd2 _7518_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7393__A _7436_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_31_244 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7449_ hold212/X _7805_/D _7451_/S vssd2 vssd2 vccd2 vccd2 _7449_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_255 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_31_299 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_98_233 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_86_406 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_98_277 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6214__A2 _5994_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7568__A _7613_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4225__A1 _4044_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_79_491 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_13_15 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_94_461 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4704__B _4704_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4776__A2 _5142_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_13_48 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7175__B1 _7222_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_81_199 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5816__A _5816_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_35_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_112_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_62_391 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_10_406 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_10_428 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_54_11 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_54_99 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6820_ _6820_/A _6820_/B _6820_/C vssd2 vssd2 vccd2 vccd2 _6822_/A sky130_fd_sc_hd__or3_2
XANTENNA__7197__B _7197_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4216__B2 _4162_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5413__B1 _4814_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6751_ _6685_/A _6685_/B _6683_/Y vssd2 vssd2 vccd2 vccd2 _6753_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_73_601 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_57_152 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_3963_ _7775_/Q _4050_/B vssd2 vssd2 vccd2 vccd2 _3964_/B sky130_fd_sc_hd__nand2_2
X_6682_ _6600_/A _6600_/B _6598_/Y vssd2 vssd2 vccd2 vccd2 _6684_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_45_325 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5702_ _7883_/Q _7884_/Q _5694_/X _5735_/B vssd2 vssd2 vccd2 vccd2 _5704_/B sky130_fd_sc_hd__o31a_2
X_3894_ _3894_/A _4083_/B _3993_/D _3893_/D vssd2 vssd2 vccd2 vccd2 _3895_/D sky130_fd_sc_hd__or4b_1
X_5633_ _7856_/Q _7855_/Q _7857_/Q _7858_/Q _5645_/B vssd2 vssd2 vccd2 vccd2 _5641_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_0_5_433 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5564_ _5573_/C _5573_/D vssd2 vssd2 vccd2 vccd2 _5566_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_52 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7303_ _7303_/A _7303_/B _7303_/C vssd2 vssd2 vccd2 vccd2 _7304_/A sky130_fd_sc_hd__or3_1
X_4515_ _4516_/A _4516_/B vssd2 vssd2 vccd2 vccd2 _4515_/Y sky130_fd_sc_hd__nor2_1
Xhold101 wbs_adr_i[3] vssd2 vssd2 vccd2 vccd2 input75/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 _7386_/Y vssd2 vssd2 vccd2 vccd2 _7454_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _7405_/X vssd2 vssd2 vccd2 vccd2 _7671_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 _7339_/X vssd2 vssd2 vccd2 vccd2 _7346_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5495_ _5528_/C _5526_/A _5528_/D _5463_/A vssd2 vssd2 vccd2 vccd2 _5496_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_111_463 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_111_441 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7234_ _7177_/A _7179_/B _7177_/B vssd2 vssd2 vccd2 vccd2 _7236_/B sky130_fd_sc_hd__a21bo_1
X_4446_ wire212/X _4881_/A2 _4965_/B vssd2 vssd2 vccd2 vccd2 _4448_/B sky130_fd_sc_hd__a21oi_2
Xhold167 _7412_/X vssd2 vssd2 vccd2 vccd2 _7413_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _7402_/X vssd2 vssd2 vccd2 vccd2 _7403_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 wbs_dat_i[15] vssd2 vssd2 vccd2 vccd2 input89/A sky130_fd_sc_hd__dlygate4sd3_1
X_7165_ _7166_/A _7166_/B _7166_/C vssd2 vssd2 vccd2 vccd2 _7167_/A sky130_fd_sc_hd__o21a_1
XANTENNA__6557__A _6783_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold178 _7390_/X vssd2 vssd2 vccd2 vccd2 _7391_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 hold386/X vssd2 vssd2 vccd2 vccd2 _7796_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4377_ _4656_/A _4160_/B _4376_/X _4814_/B vssd2 vssd2 vccd2 vccd2 _4377_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_95_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6116_ _6115_/B _6115_/C _6115_/A vssd2 vssd2 vccd2 vccd2 _6116_/X sky130_fd_sc_hd__o21a_1
XTAP_450 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _7143_/B _7222_/B _7294_/C _7143_/A vssd2 vssd2 vccd2 vccd2 _7098_/A sky130_fd_sc_hd__a22o_1
XTAP_461 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _5998_/A _5998_/B _5998_/C vssd2 vssd2 vccd2 vccd2 _6049_/C sky130_fd_sc_hd__a21bo_1
XTAP_1605 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_439 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1627 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_76_450 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6949_ _6949_/A _6949_/B vssd2 vssd2 vccd2 vccd2 _6950_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_64_634 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_48_174 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_36_336 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_51_306 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6132__B2 _7849_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6132__A1 _7848_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6467__A _7336_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold690 _7647_/Q vssd2 vssd2 vccd2 vccd2 hold690/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5643__B1 _5645_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_428 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_24_14 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_24_25 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4434__B _4704_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5946__A1 _7847_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_54_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_325 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_82_464 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_40_24 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_40_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_70_648 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_50_361 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5280_ _5211_/A _5213_/B _5211_/B vssd2 vssd2 vccd2 vccd2 _5281_/B sky130_fd_sc_hd__a21boi_2
X_4300_ _4301_/A _4303_/D vssd2 vssd2 vccd2 vccd2 _4360_/A sky130_fd_sc_hd__or2_1
XANTENNA__6674__A2 _7222_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5477__A3 _4800_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4231_ _4232_/A _4232_/B vssd2 vssd2 vccd2 vccd2 _4260_/B sky130_fd_sc_hd__and2_1
X_4162_ _4162_/A _4162_/B vssd2 vssd2 vccd2 vccd2 _4162_/X sky130_fd_sc_hd__and2_1
X_4093_ _4093_/A _4189_/B vssd2 vssd2 vccd2 vccd2 _4187_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_65_98 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_77_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7852_ _7854_/CLK _7852_/D _7611_/Y vssd2 vssd2 vccd2 vccd2 _7852_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_86 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4995_ _4845_/A _4845_/B _4925_/B _4994_/Y vssd2 vssd2 vccd2 vccd2 _4996_/B sky130_fd_sc_hd__a31o_4
X_7783_ _7787_/CLK _7783_/D _7542_/Y vssd2 vssd2 vccd2 vccd2 _7783_/Q sky130_fd_sc_hd__dfrtp_4
X_6803_ _7037_/A _7140_/A vssd2 vssd2 vccd2 vccd2 _6804_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_105_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6734_ _6734_/A _6734_/B vssd2 vssd2 vccd2 vccd2 _6746_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_58_494 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_18_303 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_18_325 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3946_ _4214_/B _4214_/C _7768_/Q vssd2 vssd2 vccd2 vccd2 _3947_/C sky130_fd_sc_hd__and3b_1
XFILLER_0_46_645 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_90_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6665_ _6665_/A _6665_/B vssd2 vssd2 vccd2 vccd2 _6667_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_177 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_317 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3877_ _3996_/B _4080_/D vssd2 vssd2 vccd2 vccd2 _4002_/C sky130_fd_sc_hd__nor2_2
XFILLER_0_103_205 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6596_ _6596_/A _6596_/B vssd2 vssd2 vccd2 vccd2 _6599_/A sky130_fd_sc_hd__xnor2_2
X_5616_ _7864_/Q _5616_/B vssd2 vssd2 vccd2 vccd2 _5620_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_249 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5547_ _5454_/A _5454_/B _5547_/C _5547_/D vssd2 vssd2 vccd2 vccd2 _5548_/B sky130_fd_sc_hd__and4bb_1
XANTENNA__7311__B1 _6069_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5478_ _5478_/A _5478_/B vssd2 vssd2 vccd2 vccd2 _5480_/C sky130_fd_sc_hd__xor2_1
X_7217_ _7279_/A _7217_/B vssd2 vssd2 vccd2 vccd2 _7310_/A sky130_fd_sc_hd__xor2_2
X_4429_ _4328_/A _4815_/B _3971_/Y _4428_/X _4025_/C vssd2 vssd2 vccd2 vccd2 _4429_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_111_293 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7148_ _7149_/A _7149_/B vssd2 vssd2 vccd2 vccd2 _7191_/A sky130_fd_sc_hd__and2b_1
X_7079_ _7081_/A _7081_/B _7081_/C vssd2 vssd2 vccd2 vccd2 _7082_/A sky130_fd_sc_hd__o21a_1
XTAP_291 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4428__B2 _4454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1424 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XTAP_1402 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5928__A1 _6670_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1479 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3939__B1 _4050_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_107_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_91_261 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_24_306 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_317 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5366__A _5366_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_10_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_10_16 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_339 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_36_188 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_51_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_20_523 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6197__A _6550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_19_36 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_87_501 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_35_46 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_35_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__6363__C _7099_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4445__A _5029_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_35_68 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_87_578 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_87_567 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_59_258 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4780_ _4780_/A _4780_/B vssd2 vssd2 vccd2 vccd2 _4789_/A sky130_fd_sc_hd__xor2_4
XANTENNA__6041__B1 _5992_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_51_23 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3800_ _6253_/A vssd2 vssd2 vccd2 vccd2 _6587_/A sky130_fd_sc_hd__inv_2
XFILLER_0_7_517 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_55_486 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_177 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5276__A _5276_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_113_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6450_ _6450_/A _6450_/B vssd2 vssd2 vccd2 vccd2 _6452_/A sky130_fd_sc_hd__xnor2_2
X_6381_ _6381_/A _6381_/B vssd2 vssd2 vccd2 vccd2 _6384_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_70_456 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5401_ _5401_/A _5401_/B vssd2 vssd2 vccd2 vccd2 _5547_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_30_309 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_11_534 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_11_523 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5332_ _5333_/A _5333_/B vssd2 vssd2 vccd2 vccd2 _5412_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_50_191 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_76_42 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5263_ _4327_/X _4331_/X _4814_/Y _4267_/D vssd2 vssd2 vccd2 vccd2 _5266_/A sky130_fd_sc_hd__o211a_1
XANTENNA__4658__A1 _4809_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5194_ _5195_/A _5195_/B vssd2 vssd2 vccd2 vccd2 _5194_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_76_75 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_76_64 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4214_ _4814_/A _4214_/B _4214_/C vssd2 vssd2 vccd2 vccd2 _4214_/Y sky130_fd_sc_hd__nor3_1
X_7002_ _7003_/A _7003_/B vssd2 vssd2 vccd2 vccd2 _7002_/X sky130_fd_sc_hd__and2b_1
X_4145_ _4143_/Y _4144_/X _4148_/C vssd2 vssd2 vccd2 vccd2 _4145_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_92_41 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6280__B1 _7140_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4076_ _7766_/Q _4458_/D _4002_/A _7764_/Q _4454_/B vssd2 vssd2 vccd2 vccd2 _4076_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_92_85 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7835_ _7838_/CLK _7835_/D _7594_/Y vssd2 vssd2 vccd2 vccd2 _7835_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4978_ _4978_/A _4978_/B vssd2 vssd2 vccd2 vccd2 _4981_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_58_291 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7766_ _7798_/CLK _7766_/D _7525_/Y vssd2 vssd2 vccd2 vccd2 _7766_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_144 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7385__B _7385_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_73_261 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6717_ _6718_/A _6718_/B vssd2 vssd2 vccd2 vccd2 _6717_/Y sky130_fd_sc_hd__nor2_1
X_7697_ _7798_/CLK _7697_/D vssd2 vssd2 vccd2 vccd2 _7697_/Q sky130_fd_sc_hd__dfxtp_1
X_3929_ _3919_/X _3920_/Y _4252_/D vssd2 vssd2 vccd2 vccd2 _3929_/Y sky130_fd_sc_hd__a21oi_1
X_6648_ _6648_/A _6648_/B vssd2 vssd2 vccd2 vccd2 _6650_/B sky130_fd_sc_hd__xor2_1
XANTENNA__4090__A _4598_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_hold104_A _7454_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_33_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6579_ _6425_/A _6430_/B _7099_/B _5931_/C vssd2 vssd2 vccd2 vccd2 _6582_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_41_180 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6638__A2 _5993_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout230 hold104/X vssd2 vssd2 vccd2 vccd2 _7485_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout263 _7850_/Q vssd2 vssd2 vccd2 vccd2 _6282_/A sky130_fd_sc_hd__buf_4
Xfanout252 hold404/X vssd2 vssd2 vccd2 vccd2 _5455_/A sky130_fd_sc_hd__clkbuf_8
Xfanout274 _7770_/Q vssd2 vssd2 vccd2 vccd2 _4162_/A sky130_fd_sc_hd__buf_4
Xfanout285 _7564_/A vssd2 vssd2 vccd2 vccd2 _7565_/A sky130_fd_sc_hd__buf_8
XFILLER_0_88_309 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1232 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6480__A _6707_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1265 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_261 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__5096__A _5220_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_92_592 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_52_412 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_107_385 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_12_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_52_489 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_110_528 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_103_591 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6655__A _6973_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5950_ _5907_/D _6634_/B _5948_/X _6436_/A vssd2 vssd2 vccd2 vccd2 _5952_/B sky130_fd_sc_hd__a22o_1
XANTENNA__6801__A2 _6430_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4901_ _4819_/A _4819_/B _4817_/X vssd2 vssd2 vccd2 vccd2 _4903_/B sky130_fd_sc_hd__a21oi_2
X_5881_ _6397_/A _6019_/D _5979_/D _5920_/D vssd2 vssd2 vccd2 vccd2 _5886_/D sky130_fd_sc_hd__and4_1
X_7620_ _7645_/A vssd2 vssd2 vccd2 vccd2 _7620_/Y sky130_fd_sc_hd__inv_2
X_4832_ _4833_/A _4833_/B vssd2 vssd2 vccd2 vccd2 _4832_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_28_442 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_90_529 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4763_ _4679_/A _4679_/B _4680_/Y vssd2 vssd2 vccd2 vccd2 _4765_/B sky130_fd_sc_hd__o21a_1
X_7551_ _7557_/A vssd2 vssd2 vccd2 vccd2 _7551_/Y sky130_fd_sc_hd__inv_2
X_6502_ _6502_/A _6502_/B vssd2 vssd2 vccd2 vccd2 _6524_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_83_592 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_55_294 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_43_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7482_ _7722_/Q _7483_/A2 _7483_/B1 hold353/X vssd2 vssd2 vccd2 vccd2 _7482_/X sky130_fd_sc_hd__a22o_1
X_4694_ _4621_/A _4621_/B _4693_/A _4556_/B _4556_/A vssd2 vssd2 vccd2 vccd2 _4849_/C
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_0_70_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_70_242 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4341__C _5030_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_43_478 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_15_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6433_ _6253_/A _5713_/Y _5752_/Y _6510_/A _6432_/X vssd2 vssd2 vccd2 vccd2 _7222_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_102_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_70_275 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4879__A1 _4810_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_43_489 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__7425__S _7451_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_30_117 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6364_ _6364_/A _6364_/B vssd2 vssd2 vccd2 vccd2 _6365_/B sky130_fd_sc_hd__xnor2_2
X_6295_ _6295_/A _6295_/B vssd2 vssd2 vccd2 vccd2 _6298_/A sky130_fd_sc_hd__xnor2_2
X_5315_ _5404_/A _5315_/B _5498_/A _5468_/A vssd2 vssd2 vccd2 vccd2 _5316_/B sky130_fd_sc_hd__or4_1
X_5246_ _5248_/A _5248_/B vssd2 vssd2 vccd2 vccd2 _5247_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_53_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7293__A2 _7255_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold16 hold16/A vssd2 vssd2 vccd2 vccd2 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd2 vssd2 vccd2 vccd2 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A vssd2 vssd2 vccd2 vccd2 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ _5178_/A _5178_/B _5178_/C vssd2 vssd2 vccd2 vccd2 _5233_/A sky130_fd_sc_hd__o21a_1
Xhold49 hold49/A vssd2 vssd2 vccd2 vccd2 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
X_4128_ _7768_/Q _4160_/B _4025_/C _4025_/D _4127_/X vssd2 vssd2 vccd2 vccd2 _4128_/X
+ sky130_fd_sc_hd__a221o_1
X_4059_ _4706_/A1 _3943_/X _4018_/X _4160_/B _7767_/Q vssd2 vssd2 vccd2 vccd2 _4059_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_66_515 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7818_ _7826_/CLK _7818_/D _7577_/Y vssd2 vssd2 vccd2 vccd2 _7818_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4813__A _5042_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_46_261 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7749_ _7750_/CLK _7749_/D _7508_/Y vssd2 vssd2 vccd2 vccd2 _7749_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_464 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_46_283 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_34_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_104_333 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_6_391 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5531__A2 _5498_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6475__A _6550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_107_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_69_397 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_526 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1073 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_548 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_72_529 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1095 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_562 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_52_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_107_193 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_80_584 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
Xhold508 la_data_in[47] vssd2 vssd2 vccd2 vccd2 hold39/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_275 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xmax_cap205 _4207_/Y vssd2 vssd2 vccd2 vccd2 _5168_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_415 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
Xhold519 hold38/X vssd2 vssd2 vccd2 vccd2 _7839_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5357__D_N _5257_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xmax_cap238 _4021_/D vssd2 vssd2 vccd2 vccd2 _4122_/D sky130_fd_sc_hd__clkbuf_2
XTAP_835 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _5100_/A _5100_/B vssd2 vssd2 vccd2 vccd2 _5101_/B sky130_fd_sc_hd__xnor2_1
XTAP_802 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6080_ _6073_/Y _6078_/Y _5664_/C vssd2 vssd2 vccd2 vccd2 _6973_/B sky130_fd_sc_hd__a21o_4
X_5031_ _5030_/A _5030_/B _5030_/C _5030_/D vssd2 vssd2 vccd2 vccd2 _5033_/C sky130_fd_sc_hd__a31oi_2
XTAP_868 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3802__A _6283_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_79_128 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_73_32 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6982_ _6982_/A _6982_/B vssd2 vssd2 vccd2 vccd2 _7005_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_109 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5933_ _6008_/A _5933_/B vssd2 vssd2 vccd2 vccd2 _5958_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4797__B1 _5528_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5864_ _5865_/A _5868_/C vssd2 vssd2 vccd2 vccd2 _5917_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_367 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_63_529 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7603_ _7627_/A vssd2 vssd2 vccd2 vccd2 _7603_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4815_ _4893_/A _4815_/B vssd2 vssd2 vccd2 vccd2 _5528_/B sky130_fd_sc_hd__nand2_8
XFILLER_0_90_348 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7534_ _7557_/A vssd2 vssd2 vccd2 vccd2 _7534_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_261 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5795_ _7846_/Q _6194_/C _6130_/C vssd2 vssd2 vccd2 vccd2 _5798_/C sky130_fd_sc_hd__and3_1
XFILLER_0_113_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4746_ _4810_/A _5528_/A vssd2 vssd2 vccd2 vccd2 _4748_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_43_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA_fanout224_A _4460_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4677_ _4677_/A _4677_/B vssd2 vssd2 vccd2 vccd2 _4679_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_264 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7465_ _7705_/Q _7454_/C _7485_/B1 hold229/X vssd2 vssd2 vccd2 vccd2 _7465_/X sky130_fd_sc_hd__a22o_1
X_6416_ _6939_/A _6973_/A _6989_/A _6973_/B vssd2 vssd2 vccd2 vccd2 _6417_/B sky130_fd_sc_hd__or4_2
XANTENNA__6279__B _7094_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7396_ hold180/X _7779_/D _7418_/S vssd2 vssd2 vccd2 vccd2 _7396_/X sky130_fd_sc_hd__mux2_1
X_6347_ _6347_/A _6347_/B vssd2 vssd2 vccd2 vccd2 _6348_/B sky130_fd_sc_hd__xor2_2
X_6278_ _6278_/A _6278_/B vssd2 vssd2 vccd2 vccd2 _6295_/A sky130_fd_sc_hd__or2_2
XANTENNA__5277__B2 _5210_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5277__A1 _5210_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5229_ _5176_/A _5174_/Y _5173_/X vssd2 vssd2 vccd2 vccd2 _5231_/B sky130_fd_sc_hd__a21o_1
XANTENNA__6777__A1 _6707_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_94_654 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XPHY_134 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_123 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_112 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_101 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_156 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_145 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_66_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_54_529 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_178 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4729__C_N _5030_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_22_426 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_34_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5374__A _5431_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_104_141 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6701__A1 _6402_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5504__A2 _5431_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_27_25 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XPHY_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_85_643 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4453__A _4898_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_57_334 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_85_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_84_175 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4600_ _4708_/A _5374_/B _4601_/B vssd2 vssd2 vccd2 vccd2 _4669_/A sky130_fd_sc_hd__or3b_1
XANTENNA__4172__B _5030_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_111_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5580_ _7863_/Q _7864_/Q _7865_/Q _7866_/Q vssd2 vssd2 vccd2 vccd2 _5581_/D sky130_fd_sc_hd__or4_1
X_4531_ _4532_/A _4532_/B vssd2 vssd2 vccd2 vccd2 _4605_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_25_286 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold316 hold316/A vssd2 vssd2 vccd2 vccd2 la_data_out[28] sky130_fd_sc_hd__buf_12
Xhold305 hold658/X vssd2 vssd2 vccd2 vccd2 hold659/A sky130_fd_sc_hd__dlygate4sd3_1
X_7250_ _7310_/A _7219_/B _7336_/A vssd2 vssd2 vccd2 vccd2 _7251_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_392 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4462_ _4896_/A _4662_/B _5099_/A _4962_/A vssd2 vssd2 vccd2 vccd2 _4462_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_40_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6201_ _6082_/A _6571_/B _6139_/B _6140_/B _6140_/A vssd2 vssd2 vccd2 vccd2 _6212_/A
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4703__B1 _5076_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_68_32 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
Xhold349 _7755_/Q vssd2 vssd2 vccd2 vccd2 hold349/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 _7742_/Q vssd2 vssd2 vccd2 vccd2 hold327/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 _7476_/X vssd2 vssd2 vccd2 vccd2 _7716_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7181_ _7181_/A _7253_/C _7181_/C vssd2 vssd2 vccd2 vccd2 _7259_/A sky130_fd_sc_hd__or3_1
X_4393_ _4393_/A _4393_/B vssd2 vssd2 vccd2 vccd2 _4394_/B sky130_fd_sc_hd__or2_1
XFILLER_0_110_177 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_610 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6132_ _7848_/Q _7313_/A _6398_/B _7849_/Q vssd2 vssd2 vccd2 vccd2 _6132_/X sky130_fd_sc_hd__a22o_1
X_6063_ _6064_/A _6064_/B vssd2 vssd2 vccd2 vccd2 _6065_/B sky130_fd_sc_hd__nor2_1
XTAP_654 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5014_ _5210_/A _5210_/B _5414_/A _5081_/C vssd2 vssd2 vccd2 vccd2 _5015_/B sky130_fd_sc_hd__or4_1
XTAP_687 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_97 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA_fanout174_A _4779_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6965_ _6967_/A _6967_/B vssd2 vssd2 vccd2 vccd2 _6965_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_610 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_88_492 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_76_643 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5916_ _5917_/A _5967_/B vssd2 vssd2 vccd2 vccd2 _5965_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_91_602 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6896_ _6896_/A _6896_/B vssd2 vssd2 vccd2 vccd2 _6897_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_48_356 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_75_186 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_75_175 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_63_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5847_ _6282_/A _5992_/B _5723_/Y _6157_/A _5944_/B vssd2 vssd2 vccd2 vccd2 _5855_/C
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_581 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5778_ _5713_/Y _5776_/Y _5777_/X vssd2 vssd2 vccd2 vccd2 _5778_/X sky130_fd_sc_hd__o21ba_2
XFILLER_0_90_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4729_ _4729_/A _5222_/A _5030_/B vssd2 vssd2 vccd2 vccd2 _4730_/B sky130_fd_sc_hd__or3b_2
XANTENNA__4810__B _5498_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7517_ _7564_/A vssd2 vssd2 vccd2 vccd2 _7517_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_264 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_114_461 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7448_ _7450_/A _7448_/B vssd2 vssd2 vccd2 vccd2 _7692_/D sky130_fd_sc_hd__and2_1
XFILLER_0_31_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_101_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7379_ hold194/X _7772_/D _7383_/S vssd2 vssd2 vccd2 vccd2 _7379_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5922__A _6282_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4170__B2 _7767_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_98_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_98_289 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4273__A _4962_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4225__A2 _4044_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_104_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4704__C _5142_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_67_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_13_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_345 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_378 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_94_495 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7175__A1 _7222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7175__B2 _7099_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_54_348 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5816__B _5816_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_105_461 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_50_543 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7478__A2 _7483_/A2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_50_554 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_10_418 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_38_79 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_89_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6663__A _6812_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6750_ _6750_/A _6750_/B vssd2 vssd2 vccd2 vccd2 _6753_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_120 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5413__B2 _4800_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3962_ _7777_/Q _3962_/B vssd2 vssd2 vccd2 vccd2 _3965_/A sky130_fd_sc_hd__xnor2_4
X_5701_ _7883_/Q _7884_/Q vssd2 vssd2 vccd2 vccd2 _5705_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_18_518 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6681_ _6681_/A _6681_/B vssd2 vssd2 vccd2 vccd2 _6684_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_55 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_3893_ _3894_/A _3893_/B _4083_/B _3893_/D vssd2 vssd2 vccd2 vccd2 _3902_/C sky130_fd_sc_hd__or4_1
XFILLER_0_70_88 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5632_ _7861_/Q _5632_/B vssd2 vssd2 vccd2 vccd2 _5811_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_60_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5563_ _5573_/C _5573_/D vssd2 vssd2 vccd2 vccd2 _5570_/B sky130_fd_sc_hd__nor2_1
X_4514_ _4514_/A _4514_/B vssd2 vssd2 vccd2 vccd2 _4516_/B sky130_fd_sc_hd__xnor2_2
X_7302_ _7302_/A _7302_/B vssd2 vssd2 vccd2 vccd2 _7303_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__7469__A2 _7483_/A2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_13_234 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_79_86 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold124 hold390/X vssd2 vssd2 vccd2 vccd2 _7767_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 input75/X vssd2 vssd2 vccd2 vccd2 _7349_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 hold674/X vssd2 vssd2 vccd2 vccd2 _7385_/B sky130_fd_sc_hd__clkbuf_2
Xhold113 _7387_/X vssd2 vssd2 vccd2 vccd2 _7418_/S sky130_fd_sc_hd__buf_6
XFILLER_0_13_256 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5494_ _5528_/C _5526_/A _5528_/D vssd2 vssd2 vccd2 vccd2 _5496_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_554 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_110_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7233_ _7264_/A _7233_/B vssd2 vssd2 vccd2 vccd2 _7239_/A sky130_fd_sc_hd__and2_1
X_4445_ _5029_/A _5042_/B vssd2 vssd2 vccd2 vccd2 _4448_/A sky130_fd_sc_hd__nor2_2
Xhold146 input89/X vssd2 vssd2 vccd2 vccd2 hold146/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 wbs_dat_i[12] vssd2 vssd2 vccd2 vccd2 input86/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 wbs_dat_i[6] vssd2 vssd2 vccd2 vccd2 input95/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7433__S _7451_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_111_475 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7164_ _7164_/A _7164_/B vssd2 vssd2 vccd2 vccd2 _7166_/C sky130_fd_sc_hd__xor2_1
Xhold179 wbs_dat_i[4] vssd2 vssd2 vccd2 vccd2 input93/A sky130_fd_sc_hd__dlygate4sd3_1
X_4376_ _4328_/A _4707_/A _3928_/X _7770_/Q vssd2 vssd2 vccd2 vccd2 _4376_/X sky130_fd_sc_hd__a22o_1
X_6115_ _6115_/A _6115_/B _6115_/C vssd2 vssd2 vccd2 vccd2 _6115_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__6557__B _7181_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_0_194 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_440 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout291_A _7629_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7095_ _7095_/A _7095_/B vssd2 vssd2 vccd2 vccd2 _7104_/A sky130_fd_sc_hd__xnor2_1
XTAP_462 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _6045_/B _6045_/C _6045_/A vssd2 vssd2 vccd2 vccd2 _6049_/B sky130_fd_sc_hd__a21o_1
XTAP_495 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_237 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6948_ _6949_/A _6949_/B vssd2 vssd2 vccd2 vccd2 _6948_/X sky130_fd_sc_hd__and2_1
XFILLER_0_76_473 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_48_186 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__3966__A1 _7772_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3966__B2 _4809_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6879_ _6973_/A _6973_/B _7224_/A _7291_/A vssd2 vssd2 vccd2 vccd2 _6919_/A sky130_fd_sc_hd__or4_1
XFILLER_0_48_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_51_318 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_17_584 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_44_381 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold680 _7668_/Q vssd2 vssd2 vccd2 vccd2 hold680/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold691 _7677_/Q vssd2 vssd2 vccd2 vccd2 hold691/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4268__A _4268_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5099__A _5099_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_24_48 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_67_462 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4434__C _4711_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5946__A2 _6281_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_82_421 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_67_484 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_27_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_40_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_35_381 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_50_340 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4382__B2 _5458_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_49_78 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4230_ _4230_/A _4230_/B vssd2 vssd2 vccd2 vccd2 _4232_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__5882__A1 _7849_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4161_ _4374_/A _4252_/C vssd2 vssd2 vccd2 vccd2 _4161_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_65_11 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_65_66 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_65_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4092_ _4134_/A _4092_/B vssd2 vssd2 vccd2 vccd2 _4189_/B sky130_fd_sc_hd__or2_2
XFILLER_0_77_204 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7851_ _7854_/CLK _7851_/D _7610_/Y vssd2 vssd2 vccd2 vccd2 _7851_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_43 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6802_ _6973_/A _6973_/B _7237_/A _7224_/A vssd2 vssd2 vccd2 vccd2 _6876_/A sky130_fd_sc_hd__or4_1
XFILLER_0_77_259 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4994_ _4842_/A _4922_/X _4924_/B vssd2 vssd2 vccd2 vccd2 _4994_/Y sky130_fd_sc_hd__a21oi_1
X_7782_ _7782_/CLK _7782_/D _7541_/Y vssd2 vssd2 vccd2 vccd2 _7782_/Q sky130_fd_sc_hd__dfrtp_4
X_6733_ _6733_/A _6733_/B vssd2 vssd2 vccd2 vccd2 _6734_/B sky130_fd_sc_hd__xor2_2
X_3945_ _4214_/C vssd2 vssd2 vccd2 vccd2 _3945_/Y sky130_fd_sc_hd__inv_2
X_6664_ _6664_/A _7099_/B _6665_/B vssd2 vssd2 vccd2 vccd2 _6664_/X sky130_fd_sc_hd__and3_1
XANTENNA__5737__A _6152_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_61_605 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_45_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_5_220 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5615_ _7864_/Q _5616_/B vssd2 vssd2 vccd2 vccd2 _5630_/B sky130_fd_sc_hd__xor2_4
X_3876_ _4458_/D _4144_/C _4326_/C _4267_/D vssd2 vssd2 vccd2 vccd2 _4148_/D sky130_fd_sc_hd__or4_1
XFILLER_0_83_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6595_ _6595_/A _6595_/B vssd2 vssd2 vccd2 vccd2 _6596_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_33_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_103_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_60_148 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5546_ _5544_/B _5523_/B _5456_/A _5490_/A _5490_/B vssd2 vssd2 vccd2 vccd2 _5547_/D
+ sky130_fd_sc_hd__a2111oi_1
XANTENNA__4373__A1 _4268_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5477_ _4893_/A _4856_/B _4800_/C _5476_/Y vssd2 vssd2 vccd2 vccd2 _5478_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_111_261 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7216_ _7216_/A _7216_/B _7216_/C vssd2 vssd2 vccd2 vccd2 _7217_/B sky130_fd_sc_hd__nand3_2
X_4428_ _4706_/A1 _4125_/B _3931_/Y _4253_/B _4454_/A vssd2 vssd2 vccd2 vccd2 _4428_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6287__B _6430_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7147_ _7100_/A _7100_/B _7098_/B vssd2 vssd2 vccd2 vccd2 _7149_/B sky130_fd_sc_hd__o21ai_1
X_4359_ _4360_/A _4360_/B _4360_/C vssd2 vssd2 vccd2 vccd2 _4420_/A sky130_fd_sc_hd__a21o_1
X_7078_ _7125_/B _7078_/B vssd2 vssd2 vccd2 vccd2 _7081_/C sky130_fd_sc_hd__nor2_1
XTAP_292 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6029_ _6029_/A _6029_/B vssd2 vssd2 vccd2 vccd2 _6032_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__7399__A _7440_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7870_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_502 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1414 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_568 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_68_248 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XTAP_1469 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_112 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_36_145 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_91_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_64_487 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_52_627 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_9_581 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5366__B _5498_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6197__B _6479_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_99_362 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_87_513 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4445__B _5042_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_248 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_74_218 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6041__A1 _6039_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_95_590 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4461__A _4810_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5276__B _5468_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_498 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5707__D _6670_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_42_126 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6380_ _6380_/A _6380_/B vssd2 vssd2 vccd2 vccd2 _6381_/B sky130_fd_sc_hd__xor2_2
X_5400_ _5445_/A _5356_/B _5352_/X vssd2 vssd2 vccd2 vccd2 _5401_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_113_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5331_ _5267_/A _5267_/B _5265_/Y vssd2 vssd2 vccd2 vccd2 _5333_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_11_513 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_100_209 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_11_546 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7001_ _7001_/A _7001_/B vssd2 vssd2 vccd2 vccd2 _7003_/B sky130_fd_sc_hd__xnor2_1
X_5262_ _5325_/A _5528_/A vssd2 vssd2 vccd2 vccd2 _5267_/A sky130_fd_sc_hd__or2_1
X_5193_ _5195_/A _5195_/B vssd2 vssd2 vccd2 vccd2 _5249_/D sky130_fd_sc_hd__nand2_1
X_4213_ _4656_/A _4020_/X _4057_/X _4454_/A vssd2 vssd2 vccd2 vccd2 _4213_/X sky130_fd_sc_hd__a22o_1
X_4144_ _4490_/A _4458_/D _4144_/C _4144_/D vssd2 vssd2 vccd2 vccd2 _4144_/X sky130_fd_sc_hd__or4_1
XFILLER_0_92_53 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_78_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6280__A1 _5816_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4075_ _7767_/Q _4075_/B vssd2 vssd2 vccd2 vccd2 _4075_/X sky130_fd_sc_hd__and2_1
XFILLER_0_92_97 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7834_ _7838_/CLK _7834_/D _7593_/Y vssd2 vssd2 vccd2 vccd2 _7834_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_65_218 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7765_ _7779_/CLK _7765_/D _7524_/Y vssd2 vssd2 vccd2 vccd2 _7765_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_309 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4977_ _4977_/A _4977_/B vssd2 vssd2 vccd2 vccd2 _4978_/B sky130_fd_sc_hd__xor2_4
X_6716_ _6718_/A _6718_/B vssd2 vssd2 vccd2 vccd2 _6716_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_46_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4594__A1 _7772_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_46_465 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7696_ _7776_/CLK _7696_/D vssd2 vssd2 vccd2 vccd2 _7696_/Q sky130_fd_sc_hd__dfxtp_1
X_3928_ _4252_/D _4063_/B vssd2 vssd2 vccd2 vccd2 _3928_/X sky130_fd_sc_hd__and2_1
XANTENNA__4594__B2 _4656_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6647_ _6647_/A _6647_/B vssd2 vssd2 vccd2 vccd2 _6648_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_73_284 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_61_435 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_413 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_46_487 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_18_178 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4090__B _4807_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3859_ _7795_/Q _3860_/B vssd2 vssd2 vccd2 vccd2 _4100_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_41_90 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6578_ _6578_/A _6578_/B vssd2 vssd2 vccd2 vccd2 _6600_/A sky130_fd_sc_hd__and2_1
XFILLER_0_14_373 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5529_ _5529_/A _5529_/B vssd2 vssd2 vccd2 vccd2 _5530_/B sky130_fd_sc_hd__nand2_1
Xfanout220 _5414_/B vssd2 vssd2 vccd2 vccd2 _5374_/B sky130_fd_sc_hd__buf_4
XANTENNA__5930__A _6664_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout264 _7849_/Q vssd2 vssd2 vccd2 vccd2 _6158_/A sky130_fd_sc_hd__buf_4
Xfanout253 _7886_/Q vssd2 vssd2 vccd2 vccd2 _5735_/B sky130_fd_sc_hd__clkbuf_8
Xfanout286 _7629_/A vssd2 vssd2 vccd2 vccd2 _7564_/A sky130_fd_sc_hd__clkbuf_8
Xfanout275 _7769_/Q vssd2 vssd2 vccd2 vccd2 _4328_/A sky130_fd_sc_hd__buf_4
XFILLER_0_96_321 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4282__B1 _4966_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6810__A3 _7313_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_96_365 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1222 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_568 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7727__RESET_B _7436_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_96_398 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1266 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_229 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__6480__B _7181_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1299 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_432 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_112_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4281__A _5042_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_21_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4585__B2 _4656_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4585__A1 _4454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_92_582 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_64_295 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5096__B _5315_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_60_490 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_103_581 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6936__A _7047_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5837__B2 _6157_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6655__B _6973_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3998__C _5458_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_99_181 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_62_45 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4900_ _4900_/A _4900_/B vssd2 vssd2 vccd2 vccd2 _4903_/A sky130_fd_sc_hd__xnor2_4
X_5880_ _7847_/Q _6253_/B _6253_/C _6191_/D vssd2 vssd2 vccd2 vccd2 _5886_/C sky130_fd_sc_hd__and4_1
X_4831_ _4757_/A _4757_/B _4755_/Y vssd2 vssd2 vccd2 vccd2 _4833_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_62_67 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_75_549 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_28_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4762_ _4762_/A _4762_/B vssd2 vssd2 vccd2 vccd2 _4765_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_262 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7550_ _7557_/A vssd2 vssd2 vccd2 vccd2 _7550_/Y sky130_fd_sc_hd__inv_2
X_6501_ _6499_/X _6501_/B vssd2 vssd2 vccd2 vccd2 _6502_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_70_221 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4693_ _4693_/A _4693_/B vssd2 vssd2 vccd2 vccd2 _7739_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_7_359 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7481_ _7721_/Q _7483_/A2 _7483_/B1 hold345/X vssd2 vssd2 vccd2 vccd2 _7481_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_3_521 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6432_ _6093_/A _6587_/B _6094_/B vssd2 vssd2 vccd2 vccd2 _6432_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_3_543 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6363_ _6590_/A _6364_/A _7099_/B vssd2 vssd2 vccd2 vccd2 _6363_/X sky130_fd_sc_hd__and3_1
XFILLER_0_11_332 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6294_ _6294_/A _6294_/B vssd2 vssd2 vccd2 vccd2 _6295_/B sky130_fd_sc_hd__xor2_1
X_5314_ _5315_/B _5498_/A _5468_/A _5404_/A vssd2 vssd2 vccd2 vccd2 _5316_/A sky130_fd_sc_hd__o22ai_1
X_5245_ _5248_/B _5248_/A vssd2 vssd2 vccd2 vccd2 _5247_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_46_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold17 hold17/A vssd2 vssd2 vccd2 vccd2 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7441__S _7451_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold28 hold28/A vssd2 vssd2 vccd2 vccd2 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A vssd2 vssd2 vccd2 vccd2 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
X_5176_ _5176_/A _5176_/B vssd2 vssd2 vccd2 vccd2 _5178_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__4366__A _4898_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4127_ _7763_/Q _4815_/B _4019_/Y _7764_/Q vssd2 vssd2 vccd2 vccd2 _4127_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5547__A_N _5454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4058_ _4162_/A _4020_/X _4057_/X _7768_/Q vssd2 vssd2 vccd2 vccd2 _4058_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_78_332 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6581__A _6581_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_78_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_93_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7817_ _7826_/CLK _7817_/D _7576_/Y vssd2 vssd2 vccd2 vccd2 _7817_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4813__B _5374_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_108_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4567__A1 _4898_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7748_ _7750_/CLK _7748_/D _7507_/Y vssd2 vssd2 vccd2 vccd2 _7748_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_476 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_74_593 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7679_ _7793_/CLK _7679_/D vssd2 vssd2 vccd2 vccd2 _7679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5925__A _7847_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_34_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_104_345 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6492__A1 _6855_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_321 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1030 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_96_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5819__B _5819_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1074 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_379 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XTAP_1096 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_240 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_65_582 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_37_262 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_114_109 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_107_161 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_92_390 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_80_541 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_52_232 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_37_295 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold509 hold39/X vssd2 vssd2 vccd2 vccd2 input42/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_825 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5030_/A _5030_/B _5030_/C _5030_/D vssd2 vssd2 vccd2 vccd2 _5160_/A sky130_fd_sc_hd__and4_2
XTAP_858 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_869 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_11 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6981_ _6982_/B _6982_/A vssd2 vssd2 vccd2 vccd2 _6981_/X sky130_fd_sc_hd__and2b_1
X_5932_ _6636_/A _6812_/A _6812_/B _6550_/A vssd2 vssd2 vccd2 vccd2 _5933_/B sky130_fd_sc_hd__o22a_1
XFILLER_0_87_151 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__5994__B1 _5781_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5863_ _5863_/A _5863_/B vssd2 vssd2 vccd2 vccd2 _5868_/C sky130_fd_sc_hd__xor2_1
X_7602_ _7627_/A vssd2 vssd2 vccd2 vccd2 _7602_/Y sky130_fd_sc_hd__inv_2
X_5794_ _5586_/B _5584_/Y _5586_/Y _5630_/B vssd2 vssd2 vccd2 vccd2 _6130_/C sky130_fd_sc_hd__o211a_2
X_4814_ _4814_/A _4814_/B vssd2 vssd2 vccd2 vccd2 _4814_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_56_571 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4745_ _4745_/A _4745_/B vssd2 vssd2 vccd2 vccd2 _5105_/B sky130_fd_sc_hd__nand2_2
X_7533_ _7565_/A vssd2 vssd2 vccd2 vccd2 _7533_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_232 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_98_41 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4676_ _4676_/A _4676_/B vssd2 vssd2 vccd2 vccd2 _4677_/B sky130_fd_sc_hd__xnor2_1
X_7464_ _7704_/Q _7454_/C _7485_/B1 hold231/X vssd2 vssd2 vccd2 vccd2 _7464_/X sky130_fd_sc_hd__a22o_1
XANTENNA_fanout217_A _5145_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_114_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_98_85 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6415_ _6973_/A _6989_/A _6973_/B _6939_/A vssd2 vssd2 vccd2 vccd2 _6415_/X sky130_fd_sc_hd__o22a_1
X_7395_ _7440_/A _7395_/B vssd2 vssd2 vccd2 vccd2 _7666_/D sky130_fd_sc_hd__and2_1
XFILLER_0_31_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_101_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6346_ _6347_/A _6347_/B vssd2 vssd2 vccd2 vccd2 _6346_/X sky130_fd_sc_hd__and2_1
X_6277_ _6276_/B _6276_/C _6276_/A vssd2 vssd2 vccd2 vccd2 _6278_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__5277__A2 _5498_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5228_ _5164_/A _5550_/B _5272_/A _5227_/Y vssd2 vssd2 vccd2 vccd2 _5231_/A sky130_fd_sc_hd__a2bb2o_1
X_5159_ _5159_/A _5159_/B vssd2 vssd2 vccd2 vccd2 _5160_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_98_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6777__A2 _7291_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_94_611 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_39_516 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_124 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_102 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_39_538 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_39_549 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_157 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_146 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_135 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_19_240 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XPHY_179 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_168 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_19_262 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_105_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_104_153 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6701__A2 _7197_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5374__B _5374_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_104_197 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_89_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_97_471 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_69_151 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_43_36 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__4453__B _5220_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XPHY_4 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_53_541 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_104_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4530_ _4530_/A _4530_/B vssd2 vssd2 vccd2 vccd2 _4532_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_574 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold306 hold306/A vssd2 vssd2 vccd2 vccd2 la_data_out[23] sky130_fd_sc_hd__buf_12
Xhold317 hold670/X vssd2 vssd2 vccd2 vccd2 hold671/A sky130_fd_sc_hd__dlygate4sd3_1
X_4461_ _4810_/A _5222_/A vssd2 vssd2 vccd2 vccd2 _4465_/A sky130_fd_sc_hd__nor2_1
X_6200_ _6307_/A _6200_/B vssd2 vssd2 vccd2 vccd2 _6242_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4703__A1 _4704_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4703__B2 _4898_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7180_ _7051_/A _7253_/D _6670_/Y _6479_/C vssd2 vssd2 vccd2 vccd2 _7181_/C sky130_fd_sc_hd__o22a_1
Xhold339 _7751_/Q vssd2 vssd2 vccd2 vccd2 hold339/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 _7470_/X vssd2 vssd2 vccd2 vccd2 _7710_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4392_ _4393_/A _4393_/B vssd2 vssd2 vccd2 vccd2 _4468_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_21_471 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_600 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _6670_/A _6253_/C _6075_/D _6017_/B _7850_/Q vssd2 vssd2 vccd2 vccd2 _6131_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_110_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_68_99 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_68_88 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__6396__A _6670_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_21_493 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_611 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6062_/A _6062_/B vssd2 vssd2 vccd2 vccd2 _6065_/A sky130_fd_sc_hd__nor2_1
XTAP_655 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_65 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5013_ _5210_/B _5414_/A _5081_/C _4711_/A vssd2 vssd2 vccd2 vccd2 _5013_/X sky130_fd_sc_hd__o22a_1
XTAP_688 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_95_408 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6964_ _6964_/A _6964_/B vssd2 vssd2 vccd2 vccd2 _6967_/B sky130_fd_sc_hd__xnor2_2
X_5915_ _5915_/A _5915_/B vssd2 vssd2 vccd2 vccd2 _5967_/B sky130_fd_sc_hd__xnor2_2
X_6895_ _6896_/A _6896_/B vssd2 vssd2 vccd2 vccd2 _6895_/X sky130_fd_sc_hd__and2_1
X_5846_ _7846_/Q _5937_/B vssd2 vssd2 vccd2 vccd2 _5846_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_198 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_8_432 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_429 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5777_ _6158_/A _5992_/B _5992_/C _5769_/X _6157_/A vssd2 vssd2 vccd2 vccd2 _5777_/X
+ sky130_fd_sc_hd__a32o_1
X_4728_ _4728_/A _4728_/B vssd2 vssd2 vccd2 vccd2 _4730_/A sky130_fd_sc_hd__xnor2_2
X_7516_ _7564_/A vssd2 vssd2 vccd2 vccd2 _7516_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_102_602 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4659_ _5468_/A vssd2 vssd2 vccd2 vccd2 _4954_/C sky130_fd_sc_hd__inv_2
X_7447_ hold194/X _7804_/D _7451_/S vssd2 vssd2 vccd2 vccd2 _7447_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_473 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7378_ _7452_/A _7378_/B vssd2 vssd2 vccd2 vccd2 _7659_/D sky130_fd_sc_hd__and2_1
XFILLER_0_101_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6329_ _6402_/A _6404_/D _6330_/C vssd2 vssd2 vccd2 vccd2 _6329_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6998__A2 _7181_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4554__A _5455_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4273__B _4896_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_39_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4630__B1 _5076_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4704__D _5076_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_109_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7175__A2 _7222_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_54_316 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_82_658 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_35_552 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_2_608 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_105_473 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_38_69 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6663__B _7291_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_54_35 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_89_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_58_611 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3961_ _7776_/Q _7775_/Q _4050_/B vssd2 vssd2 vccd2 vccd2 _3962_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_57_132 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5700_ _6283_/B _6094_/B vssd2 vssd2 vccd2 vccd2 _5700_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85_496 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6680_ _6680_/A _6680_/B vssd2 vssd2 vccd2 vccd2 _6681_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_67 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_57_176 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_57_165 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3892_ _4519_/B _3892_/B _3892_/C vssd2 vssd2 vccd2 vccd2 _3892_/X sky130_fd_sc_hd__and3_1
XFILLER_0_73_669 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_72_135 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_45_349 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5758__A_N _6152_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5631_ _6253_/B _6253_/C _6018_/D vssd2 vssd2 vccd2 vccd2 _5631_/X sky130_fd_sc_hd__and3_1
X_5562_ _5561_/A _5522_/C _5561_/C _5560_/Y _5561_/X vssd2 vssd2 vccd2 vccd2 _5573_/D
+ sky130_fd_sc_hd__o311a_1
X_4513_ _4513_/A _4513_/B vssd2 vssd2 vccd2 vccd2 _4514_/B sky130_fd_sc_hd__xnor2_2
X_7301_ _7301_/A _7301_/B vssd2 vssd2 vccd2 vccd2 _7302_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_53_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_13_202 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_13_213 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_79_65 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7232_ _7232_/A _7232_/B _7232_/C vssd2 vssd2 vccd2 vccd2 _7233_/B sky130_fd_sc_hd__nand3_1
Xhold114 _7410_/X vssd2 vssd2 vccd2 vccd2 _7411_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 _7369_/X vssd2 vssd2 vccd2 vccd2 _7370_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 _7349_/Y vssd2 vssd2 vccd2 vccd2 _7454_/A sky130_fd_sc_hd__buf_1
X_5493_ _5468_/A _5528_/B _5550_/B _5414_/B vssd2 vssd2 vccd2 vccd2 _5528_/D sky130_fd_sc_hd__o22a_1
X_4444_ _4729_/A _4966_/A _5030_/B vssd2 vssd2 vccd2 vccd2 _4449_/A sky130_fd_sc_hd__or3b_4
Xhold147 _7383_/X vssd2 vssd2 vccd2 vccd2 _7384_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _7385_/Y vssd2 vssd2 vccd2 vccd2 _7420_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 input86/X vssd2 vssd2 vccd2 vccd2 hold158/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_487 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7163_ _7045_/A _7291_/B _7162_/Y vssd2 vssd2 vccd2 vccd2 _7164_/B sky130_fd_sc_hd__o21a_1
Xhold169 input95/X vssd2 vssd2 vccd2 vccd2 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
X_4375_ _4454_/A _4030_/X _4373_/X _4125_/C _4374_/Y vssd2 vssd2 vccd2 vccd2 _4375_/X
+ sky130_fd_sc_hd__a221o_1
X_6114_ _6111_/Y _6112_/X _6048_/X _6051_/X vssd2 vssd2 vccd2 vccd2 _6115_/C sky130_fd_sc_hd__a211oi_2
X_7094_ _7094_/A _7294_/B vssd2 vssd2 vccd2 vccd2 _7095_/B sky130_fd_sc_hd__nand2_1
XTAP_430 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6045_/A _6045_/B _6045_/C vssd2 vssd2 vccd2 vccd2 _6049_/A sky130_fd_sc_hd__nand3_1
XTAP_452 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout284_A _7629_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4860__B1 _5076_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_95_205 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_68_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_249 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6947_ _6862_/A _6862_/B _6859_/X vssd2 vssd2 vccd2 vccd2 _6949_/B sky130_fd_sc_hd__o21bai_1
XFILLER_0_48_165 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_48_154 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_36_316 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6878_ _6571_/B _7099_/B _7222_/B _6571_/A vssd2 vssd2 vccd2 vccd2 _6881_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_8_262 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5829_ _7847_/Q _5608_/Y _5620_/B _5630_/B _5828_/X vssd2 vssd2 vccd2 vccd2 _5829_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_91_499 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_44_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_102_421 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_114_281 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_102_487 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold670 _7824_/Q vssd2 vssd2 vccd2 vccd2 hold670/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 _7659_/Q vssd2 vssd2 vccd2 vccd2 hold681/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 _7674_/Q vssd2 vssd2 vccd2 vccd2 hold692/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5099__B _5374_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4434__D _4782_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_82_433 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6356__B1 _7237_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_54_135 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_23_522 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_360 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5843__A _6550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6939__A _6939_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_105_281 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4160_ _7769_/Q _4160_/B vssd2 vssd2 vccd2 vccd2 _4171_/B sky130_fd_sc_hd__and2_1
X_4091_ _4598_/A _4807_/A _4090_/C vssd2 vssd2 vccd2 vccd2 _4092_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_65_78 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7850_ _7854_/CLK _7850_/D _7609_/Y vssd2 vssd2 vccd2 vccd2 _7850_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4194__A _5548_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6801_ _6571_/B _6430_/B _7099_/B _6571_/A vssd2 vssd2 vccd2 vccd2 _6804_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_105_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4993_ _4993_/A _4993_/B vssd2 vssd2 vccd2 vccd2 _5128_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_58_441 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7781_ _7782_/CLK _7781_/D _7540_/Y vssd2 vssd2 vccd2 vccd2 _7781_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_85_271 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6732_ _6733_/A _6733_/B vssd2 vssd2 vccd2 vccd2 _6732_/X sky130_fd_sc_hd__and2_1
X_3944_ _7781_/Q _3944_/B vssd2 vssd2 vccd2 vccd2 _4214_/C sky130_fd_sc_hd__xor2_4
X_6663_ _6812_/A _7291_/A vssd2 vssd2 vccd2 vccd2 _6665_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_45_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3875_ _4458_/D _4144_/C _4326_/C _4267_/D vssd2 vssd2 vccd2 vccd2 _4002_/B sky130_fd_sc_hd__nor4_4
XFILLER_0_73_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_628 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5614_ _7863_/Q _5581_/A _5581_/B _5581_/C _5645_/B vssd2 vssd2 vccd2 vccd2 _5616_/B
+ sky130_fd_sc_hd__o41a_2
X_6594_ _6595_/A _6595_/B vssd2 vssd2 vccd2 vccd2 _6594_/X sky130_fd_sc_hd__and2_1
XFILLER_0_53_190 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5545_ _5561_/C _5545_/B vssd2 vssd2 vccd2 vccd2 _5549_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_352 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_76_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5476_ _5476_/A _5476_/B vssd2 vssd2 vccd2 vccd2 _5476_/Y sky130_fd_sc_hd__xnor2_1
X_7215_ _7211_/C _7127_/X _7211_/D _7214_/Y _7171_/B vssd2 vssd2 vccd2 vccd2 _7216_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_1_460 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4427_ _4427_/A _4427_/B vssd2 vssd2 vccd2 vccd2 _4427_/X sky130_fd_sc_hd__and2_1
XFILLER_0_111_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7146_ _7146_/A _7146_/B vssd2 vssd2 vccd2 vccd2 _7149_/A sky130_fd_sc_hd__xor2_1
XTAP_260 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4358_ _4418_/B _4358_/B vssd2 vssd2 vccd2 vccd2 _4360_/C sky130_fd_sc_hd__xnor2_1
X_7077_ _7077_/A _7077_/B vssd2 vssd2 vccd2 vccd2 _7078_/B sky130_fd_sc_hd__and2_1
XTAP_293 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _4289_/A _4289_/B vssd2 vssd2 vccd2 vccd2 _4291_/B sky130_fd_sc_hd__xor2_2
X_6028_ _6812_/A _6783_/A vssd2 vssd2 vccd2 vccd2 _6029_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_96_514 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XTAP_1415 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6586__B1 _7253_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_49_430 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5389__A1 _5328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1459 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_513 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_76_293 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_49_496 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_64_499 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_17_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_32_352 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_32_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_32_385 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6494__A _6571_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_99_374 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_87_558 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6041__A2 _6040_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_433 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4461__B _5222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_113_505 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6669__A _6670_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_23_352 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_23_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5330_ _5330_/A _5330_/B vssd2 vssd2 vccd2 vccd2 _5333_/A sky130_fd_sc_hd__xnor2_2
X_5261_ _5145_/A _5431_/B _5260_/X vssd2 vssd2 vccd2 vccd2 _5297_/A sky130_fd_sc_hd__o21ai_2
X_4212_ _7768_/Q _4030_/X _4210_/X _3971_/Y _4211_/X vssd2 vssd2 vccd2 vccd2 _4212_/X
+ sky130_fd_sc_hd__a221o_1
X_7000_ _7001_/A _7001_/B vssd2 vssd2 vccd2 vccd2 _7000_/Y sky130_fd_sc_hd__nand2b_1
X_5192_ _5192_/A _5192_/B vssd2 vssd2 vccd2 vccd2 _5195_/B sky130_fd_sc_hd__xnor2_4
X_4143_ _7768_/Q _4458_/D vssd2 vssd2 vccd2 vccd2 _4143_/Y sky130_fd_sc_hd__nand2_1
X_4074_ _7768_/Q _4326_/C _3899_/D _4162_/A vssd2 vssd2 vccd2 vccd2 _4074_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6280__A2 _5816_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_92_65 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7833_ _7838_/CLK _7833_/D _7592_/Y vssd2 vssd2 vccd2 vccd2 _7833_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_558 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7764_ _7800_/CLK _7764_/D _7523_/Y vssd2 vssd2 vccd2 vccd2 _7764_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__7439__S _7451_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4976_ _4977_/A _4977_/B vssd2 vssd2 vccd2 vccd2 _4976_/Y sky130_fd_sc_hd__nor2_1
X_6715_ _6855_/A _7181_/A _6643_/A _6640_/Y vssd2 vssd2 vccd2 vccd2 _6718_/B sky130_fd_sc_hd__o31ai_2
XFILLER_0_46_433 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_46_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7695_ _7776_/CLK _7695_/D vssd2 vssd2 vccd2 vccd2 _7695_/Q sky130_fd_sc_hd__dfxtp_1
X_3927_ _3927_/A _3927_/B _4050_/B vssd2 vssd2 vccd2 vccd2 _3982_/B sky130_fd_sc_hd__nor3b_4
X_6646_ _6647_/A _6647_/B vssd2 vssd2 vccd2 vccd2 _6646_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_46_499 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_6_541 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3858_ _3858_/A _3858_/B vssd2 vssd2 vccd2 vccd2 _4080_/D sky130_fd_sc_hd__and2_2
X_6577_ _6576_/B _6576_/C _6576_/A vssd2 vssd2 vccd2 vccd2 _6578_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__6740__B1 _6669_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_61_447 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5528_ _5528_/A _5528_/B _5528_/C _5528_/D vssd2 vssd2 vccd2 vccd2 _5529_/B sky130_fd_sc_hd__or4_1
X_5459_ _5459_/A _5528_/C vssd2 vssd2 vccd2 vccd2 _5462_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4099__A _7765_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout210 _4072_/Y vssd2 vssd2 vccd2 vccd2 _4807_/A sky130_fd_sc_hd__clkbuf_4
Xfanout221 _5081_/C vssd2 vssd2 vccd2 vccd2 _5406_/A sky130_fd_sc_hd__clkbuf_8
Xfanout232 _6588_/B vssd2 vssd2 vccd2 vccd2 _6510_/B sky130_fd_sc_hd__clkbuf_8
X_7129_ _7211_/A _7128_/X _7127_/X vssd2 vssd2 vccd2 vccd2 _7130_/B sky130_fd_sc_hd__o21a_1
Xfanout254 _7870_/Q vssd2 vssd2 vccd2 vccd2 _5645_/B sky130_fd_sc_hd__clkbuf_8
Xfanout265 _7848_/Q vssd2 vssd2 vccd2 vccd2 _6157_/A sky130_fd_sc_hd__buf_4
Xfanout243 _4253_/B vssd2 vssd2 vccd2 vccd2 _4252_/D sky130_fd_sc_hd__buf_4
Xfanout287 _7629_/A vssd2 vssd2 vccd2 vccd2 _7641_/A sky130_fd_sc_hd__buf_8
Xfanout276 _7454_/C vssd2 vssd2 vccd2 vccd2 _7483_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_69_536 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4282__A1 _4044_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_96_333 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1223 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_377 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_84_517 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XTAP_1256 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4562__A _4736_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1289 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_230 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5584__B1_N _5645_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4281__B _5029_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_21_17 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_25_617 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_37_444 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_52_425 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_9_390 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_32_171 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6936__B _7222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_20_399 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6655__C _7045_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_46_58 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_99_193 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_87_344 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_4830_ _4830_/A _4830_/B vssd2 vssd2 vccd2 vccd2 _4833_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_87_366 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_62_79 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_47_208 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_28_400 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_83_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4761_ _4759_/Y _4761_/B vssd2 vssd2 vccd2 vccd2 _4762_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_55_252 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_55_241 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6500_ _6500_/A _6500_/B _6500_/C vssd2 vssd2 vccd2 vccd2 _6501_/B sky130_fd_sc_hd__or3_1
X_4692_ _4557_/B _4622_/B _5455_/A vssd2 vssd2 vccd2 vccd2 _4693_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_7_349 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7480_ _7720_/Q _7483_/A2 _7483_/B1 hold351/X vssd2 vssd2 vccd2 vccd2 _7480_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_102_41 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6431_ _5816_/A _5816_/B _7224_/A vssd2 vssd2 vccd2 vccd2 _6437_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_113_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6362_ _6590_/A _7099_/B vssd2 vssd2 vccd2 vccd2 _6364_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4879__A3 _5498_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_23_193 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5313_ _5313_/A _5313_/B vssd2 vssd2 vccd2 vccd2 _5320_/A sky130_fd_sc_hd__xnor2_1
X_6293_ _6294_/A _6294_/B vssd2 vssd2 vccd2 vccd2 _6293_/Y sky130_fd_sc_hd__nor2_1
X_5244_ _5192_/A _5190_/Y _5189_/Y vssd2 vssd2 vccd2 vccd2 _5248_/B sky130_fd_sc_hd__a21oi_1
Xhold29 hold29/A vssd2 vssd2 vccd2 vccd2 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
X_5175_ _5175_/A _5175_/B vssd2 vssd2 vccd2 vccd2 _5176_/B sky130_fd_sc_hd__xor2_1
Xhold18 hold18/A vssd2 vssd2 vccd2 vccd2 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
X_4126_ _4268_/A _4029_/X _4030_/X _7766_/Q _4125_/X vssd2 vssd2 vccd2 vccd2 _4126_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA_fanout197_A _4318_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4366__B _4863_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4057_ _4162_/B _4125_/C _4057_/C vssd2 vssd2 vccd2 vccd2 _4057_/X sky130_fd_sc_hd__and3_1
XANTENNA__6581__B _7140_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7816_ _7826_/CLK _7816_/D _7575_/Y vssd2 vssd2 vccd2 vccd2 _7816_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_208 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_38_219 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_78_399 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__4567__A2 _5276_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4959_ _4960_/B _4959_/B vssd2 vssd2 vccd2 vccd2 _5024_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_46_241 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7747_ _7771_/CLK _7747_/D _7506_/Y vssd2 vssd2 vccd2 vccd2 _7747_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_200 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7678_ _7771_/CLK _7678_/D vssd2 vssd2 vccd2 vccd2 _7678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_499 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_233 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6629_ _6670_/A _6629_/B _6629_/C vssd2 vssd2 vccd2 vccd2 _7291_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_104_357 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6102__A _6253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_30_642 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6492__A2 _6572_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6475__C _7253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4557__A _5455_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_16_17 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4255__A1 _7767_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_333 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_96_141 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_69_366 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1031 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_517 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5819__C _6402_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1064 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5204__B1 _5498_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_32_16 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1097 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_37_285 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6704__B1 _7253_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_52_266 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_597 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_103_390 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_57_35 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XTAP_826 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_558 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6666__B _7237_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_57_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XTAP_859 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_108 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6980_ _7060_/A _6979_/X _6873_/A _6670_/Y vssd2 vssd2 vccd2 vccd2 _6982_/B sky130_fd_sc_hd__o2bb2a_1
X_5931_ _6550_/A _6402_/A _5931_/C _6664_/A vssd2 vssd2 vccd2 vccd2 _6008_/A sky130_fd_sc_hd__and4b_2
XFILLER_0_73_89 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5994__A1 _5991_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5862_ _5862_/A _5862_/B vssd2 vssd2 vccd2 vccd2 _5863_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_358 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4813_ _5042_/A _5374_/B vssd2 vssd2 vccd2 vccd2 _4818_/A sky130_fd_sc_hd__or2_2
XFILLER_0_7_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7601_ _7627_/A vssd2 vssd2 vccd2 vccd2 _7601_/Y sky130_fd_sc_hd__inv_2
X_5793_ _5607_/A _5607_/B _5620_/B _5653_/C _5599_/B vssd2 vssd2 vccd2 vccd2 _6194_/C
+ sky130_fd_sc_hd__o2111a_2
XFILLER_0_113_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7532_ _7564_/A vssd2 vssd2 vccd2 vccd2 _7532_/Y sky130_fd_sc_hd__inv_2
X_4744_ _4745_/A _4745_/B vssd2 vssd2 vccd2 vccd2 _5030_/C sky130_fd_sc_hd__and2_2
XFILLER_0_98_53 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4675_ _4676_/A _4676_/B vssd2 vssd2 vccd2 vccd2 _4675_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_71_575 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7463_ _7703_/Q _7454_/C _7485_/B1 hold243/X vssd2 vssd2 vccd2 vccd2 _7463_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_16_469 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_101_305 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6414_ _6354_/A _6354_/B _6352_/X vssd2 vssd2 vccd2 vccd2 _6421_/A sky130_fd_sc_hd__a21oi_2
X_7394_ hold207/X _7666_/Q _7418_/S vssd2 vssd2 vccd2 vccd2 _7394_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_491 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6345_ _6345_/A _6345_/B vssd2 vssd2 vccd2 vccd2 _6347_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_97 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6276_ _6276_/A _6276_/B _6276_/C vssd2 vssd2 vccd2 vccd2 _6278_/A sky130_fd_sc_hd__and3_1
X_5227_ _5227_/A _5227_/B _5227_/C vssd2 vssd2 vccd2 vccd2 _5227_/Y sky130_fd_sc_hd__nand3_1
X_5158_ _5158_/A _5158_/B vssd2 vssd2 vccd2 vccd2 _5159_/B sky130_fd_sc_hd__or2_1
X_5089_ _5089_/A _5089_/B vssd2 vssd2 vccd2 vccd2 _5089_/Y sky130_fd_sc_hd__xnor2_1
X_4109_ _4490_/A _4458_/C _4141_/C _4141_/D vssd2 vssd2 vccd2 vccd2 _4109_/X sky130_fd_sc_hd__or4_1
XFILLER_0_2_70 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_78_130 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_109_405 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_93_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_78_185 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XPHY_125 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_114 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_103 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_158 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_147 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_136 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_47_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_74_380 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_62_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_104_121 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_62_586 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_62_575 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_22_439 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5374__C _5468_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_104_165 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_30_461 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7598__A _7627_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5976__A1 _7845_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5976__B2 _7846_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XPHY_5 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_84_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_38_550 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_72_306 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5846__A _7846_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_25_244 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_25_266 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold307 hold660/X vssd2 vssd2 vccd2 vccd2 hold661/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_439 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4460_ _4456_/X _4457_/X _4458_/X _4459_/Y _4006_/C vssd2 vssd2 vccd2 vccd2 _4460_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_40_214 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
Xhold318 hold318/A vssd2 vssd2 vccd2 vccd2 la_data_out[17] sky130_fd_sc_hd__buf_12
XANTENNA__4703__A2 _5142_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4391_ _4391_/A _4391_/B vssd2 vssd2 vccd2 vccd2 _4393_/B sky130_fd_sc_hd__xnor2_1
Xhold329 _7743_/Q vssd2 vssd2 vccd2 vccd2 hold329/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_67 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_68_56 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__3911__B1 _4050_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_21_483 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6130_ _6398_/A _6194_/C _6130_/C vssd2 vssd2 vccd2 vccd2 _6130_/X sky130_fd_sc_hd__and3_1
XTAP_601 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _6059_/A _6064_/B _6128_/A _6059_/D vssd2 vssd2 vccd2 vccd2 _6062_/B sky130_fd_sc_hd__o22a_1
XANTENNA__4197__A _5548_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_656 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5012_/A _5012_/B vssd2 vssd2 vccd2 vccd2 _5022_/A sky130_fd_sc_hd__xor2_2
XTAP_678 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_88_450 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6963_ _6963_/A _6963_/B vssd2 vssd2 vccd2 vccd2 _6964_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_17_93 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_76_645 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5914_ _5915_/A _5915_/B vssd2 vssd2 vccd2 vccd2 _5962_/B sky130_fd_sc_hd__nand2b_1
X_6894_ _6826_/A _6826_/B _6824_/X vssd2 vssd2 vccd2 vccd2 _6896_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_48_347 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5845_ _6154_/A _5845_/B _5845_/C _5755_/C vssd2 vssd2 vccd2 vccd2 _5845_/X sky130_fd_sc_hd__or4b_1
XANTENNA__4660__A _4810_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_8_455 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7447__S _7451_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_29_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_92 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_106_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_8_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5776_ _7843_/Q _6094_/B _5775_/Y vssd2 vssd2 vccd2 vccd2 _5776_/Y sky130_fd_sc_hd__a21boi_1
X_4727_ _4728_/A _4728_/B vssd2 vssd2 vccd2 vccd2 _4727_/Y sky130_fd_sc_hd__nand2_1
X_7515_ _7564_/A vssd2 vssd2 vccd2 vccd2 _7515_/Y sky130_fd_sc_hd__inv_2
X_7446_ _7452_/A _7446_/B vssd2 vssd2 vccd2 vccd2 _7691_/D sky130_fd_sc_hd__and2_1
XFILLER_0_16_277 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4658_ _4809_/A _4103_/B _4656_/X _4657_/X vssd2 vssd2 vccd2 vccd2 _4880_/B sky130_fd_sc_hd__o211ai_4
XFILLER_0_101_113 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xinput90 input90/A vssd2 vssd2 vccd2 vccd2 input90/X sky130_fd_sc_hd__clkbuf_1
X_4589_ _4810_/A _5406_/A vssd2 vssd2 vccd2 vccd2 _4593_/A sky130_fd_sc_hd__nor2_1
X_7377_ hold158/X _7659_/Q _7383_/S vssd2 vssd2 vccd2 vccd2 _7377_/X sky130_fd_sc_hd__mux2_1
X_6328_ _6402_/A _6404_/D _6330_/C vssd2 vssd2 vccd2 vccd2 _6331_/A sky130_fd_sc_hd__a21oi_1
X_6259_ _6259_/A _6259_/B vssd2 vssd2 vccd2 vccd2 _6261_/C sky130_fd_sc_hd__xor2_1
XANTENNA__6852__C1 _5992_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_66_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_94_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4630__A1 _4736_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4630__B2 _4708_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_66_144 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_369 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_358 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7357__S _7383_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_109_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_81_147 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_81_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_62_361 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7332__B1 _7336_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_62_383 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6497__A _6939_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4729__B _5222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_38_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_3960_ _4018_/B _4036_/B vssd2 vssd2 vccd2 vccd2 _4025_/D sky130_fd_sc_hd__and2_1
XFILLER_0_18_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_85_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3891_ _4454_/B _7763_/Q _7791_/Q vssd2 vssd2 vccd2 vccd2 _3892_/C sky130_fd_sc_hd__and3b_1
X_5630_ _6191_/D _5630_/B _6075_/C _6019_/C vssd2 vssd2 vccd2 vccd2 _6018_/D sky130_fd_sc_hd__nor4_2
X_5561_ _5561_/A _5561_/B _5561_/C vssd2 vssd2 vccd2 vccd2 _5561_/X sky130_fd_sc_hd__or3_1
X_4512_ _4513_/A _4513_/B vssd2 vssd2 vccd2 vccd2 _4512_/Y sky130_fd_sc_hd__nand2_1
X_7300_ _7300_/A _7300_/B vssd2 vssd2 vccd2 vccd2 _7301_/B sky130_fd_sc_hd__or2_1
X_5492_ _5492_/A _5492_/B vssd2 vssd2 vccd2 vccd2 _7752_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_597 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_110_41 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7231_ _7232_/A _7232_/B _7232_/C vssd2 vssd2 vccd2 vccd2 _7264_/A sky130_fd_sc_hd__a21o_1
Xhold115 _7411_/X vssd2 vssd2 vccd2 vccd2 _7674_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 wbs_dat_i[10] vssd2 vssd2 vccd2 vccd2 input84/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 _7454_/Y vssd2 vssd2 vccd2 vccd2 hold104/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_85 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_79_99 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4443_ _4810_/A _4965_/B _4388_/X _4390_/B vssd2 vssd2 vccd2 vccd2 _4451_/A sky130_fd_sc_hd__o31a_2
Xhold137 _7441_/X vssd2 vssd2 vccd2 vccd2 _7442_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 _7377_/X vssd2 vssd2 vccd2 vccd2 _7378_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 hold389/X vssd2 vssd2 vccd2 vccd2 _7806_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7162_ _7162_/A _7162_/B vssd2 vssd2 vccd2 vccd2 _7162_/Y sky130_fd_sc_hd__xnor2_1
X_4374_ _4374_/A _4814_/B vssd2 vssd2 vccd2 vccd2 _4374_/Y sky130_fd_sc_hd__nor2_1
X_6113_ _6048_/X _6051_/X _6111_/Y _6112_/X vssd2 vssd2 vccd2 vccd2 _6115_/B sky130_fd_sc_hd__o211a_1
X_7093_ _7093_/A _7093_/B vssd2 vssd2 vccd2 vccd2 _7095_/A sky130_fd_sc_hd__nand2_1
XTAP_420 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _6105_/A _6105_/B _6939_/A _6989_/A vssd2 vssd2 vccd2 vccd2 _6045_/C sky130_fd_sc_hd__or4_1
XTAP_453 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_70 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_28_92 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4860__A1 _5168_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_fanout277_A _7453_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4860__B2 _4704_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1619 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6946_ _6946_/A _6946_/B vssd2 vssd2 vccd2 vccd2 _6949_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_442 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_91_401 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_64_604 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6877_ _6815_/A _6815_/C _6811_/X vssd2 vssd2 vccd2 vccd2 _6883_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_36_306 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5828_ _7845_/Q _5828_/B _5828_/C vssd2 vssd2 vccd2 vccd2 _5828_/X sky130_fd_sc_hd__and3_1
XFILLER_0_91_478 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_63_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_63_147 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5759_ _6152_/C _6281_/C _5759_/C vssd2 vssd2 vccd2 vccd2 _5760_/D sky130_fd_sc_hd__and3_1
XFILLER_0_44_372 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_44_361 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_17_575 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_411 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_32_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_114_293 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_102_433 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7429_ hold180/X _7795_/D _7451_/S vssd2 vssd2 vccd2 vccd2 _7429_/X sky130_fd_sc_hd__mux2_1
Xhold660 _7838_/Q vssd2 vssd2 vccd2 vccd2 hold660/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_102_455 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold671 hold671/A vssd2 vssd2 vccd2 vccd2 hold671/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 _7658_/Q vssd2 vssd2 vccd2 vccd2 hold693/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 _7671_/Q vssd2 vssd2 vccd2 vccd2 hold682/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_17 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_67_420 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_39_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_55_615 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_54_103 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_306 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6356__A1 _5816_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_70_607 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_42_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_40_49 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__5843__B _6092_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_62_191 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6939__B _7255_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_105_293 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_65_46 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4090_ _4598_/A _4807_/A _4090_/C vssd2 vssd2 vccd2 vccd2 _4134_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_77_239 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6800_ _6737_/A _6739_/B _6737_/B vssd2 vssd2 vccd2 vccd2 _6806_/A sky130_fd_sc_hd__o21bai_1
X_4992_ _4993_/A _4993_/B vssd2 vssd2 vccd2 vccd2 _4992_/Y sky130_fd_sc_hd__nor2_1
X_7780_ _7782_/CLK _7780_/D _7539_/Y vssd2 vssd2 vccd2 vccd2 _7780_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_92_209 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6731_ _6731_/A _6731_/B vssd2 vssd2 vccd2 vccd2 _6733_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_486 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_3943_ _4315_/B _4427_/A vssd2 vssd2 vccd2 vccd2 _3943_/X sky130_fd_sc_hd__and2_1
X_6662_ _6664_/A _7099_/B vssd2 vssd2 vccd2 vccd2 _6665_/A sky130_fd_sc_hd__nand2_1
X_3874_ _3813_/A _3813_/B _4745_/A _4454_/B _4656_/C vssd2 vssd2 vccd2 vccd2 _4148_/C
+ sky130_fd_sc_hd__a2111o_2
XFILLER_0_73_467 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_45_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_45_158 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5613_ _5581_/A _5581_/B _5581_/C _5645_/B vssd2 vssd2 vccd2 vccd2 _5619_/B sky130_fd_sc_hd__o31a_2
XFILLER_0_73_489 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6593_ _6668_/A _7099_/B _6516_/B _6514_/X vssd2 vssd2 vccd2 vccd2 _6595_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_14_512 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_60_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5544_ _5516_/A _5544_/B vssd2 vssd2 vccd2 vccd2 _5545_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_30_82 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_30_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5475_ _5475_/A _5475_/B _5476_/B vssd2 vssd2 vccd2 vccd2 _5512_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_41_364 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7214_ _7126_/A _7214_/B vssd2 vssd2 vccd2 vccd2 _7214_/Y sky130_fd_sc_hd__nand2b_1
X_4426_ _4162_/A _4707_/A _4063_/X _7772_/Q vssd2 vssd2 vccd2 vccd2 _4427_/B sky130_fd_sc_hd__a22o_1
X_7145_ _7145_/A _7222_/B vssd2 vssd2 vccd2 vccd2 _7146_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_472 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_250 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4357_ _4299_/A _4299_/B _4296_/X vssd2 vssd2 vccd2 vccd2 _4358_/B sky130_fd_sc_hd__a21oi_1
X_7076_ _7077_/A _7077_/B vssd2 vssd2 vccd2 vccd2 _7125_/B sky130_fd_sc_hd__nor2_1
X_4288_ _4289_/A _4289_/B vssd2 vssd2 vccd2 vccd2 _4323_/B sky130_fd_sc_hd__and2_1
XTAP_261 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6027_ _6138_/A _6812_/B vssd2 vssd2 vccd2 vccd2 _6029_/A sky130_fd_sc_hd__nor2_1
XTAP_294 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6586__A1 _5816_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_49_442 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5389__A2 _5431_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1449 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_464 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_49_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6929_ _6930_/A _6930_/B vssd2 vssd2 vccd2 vccd2 _6982_/A sky130_fd_sc_hd__and2_1
XANTENNA__6338__A1 _6634_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_64_434 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_24_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_107_569 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_45_670 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5944__A _6282_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_44_180 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_32_342 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
Xhold490 input7/X vssd2 vssd2 vccd2 vccd2 hold28/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_386 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_87_537 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6329__A1 _6402_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_82_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_55_478 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_55_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_27_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_70_437 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_70_404 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_113_517 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6669__B _6670_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5260_ _5260_/A _5260_/B vssd2 vssd2 vccd2 vccd2 _5260_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_23_397 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4211_ _7765_/Q _4815_/B _4019_/Y _7766_/Q vssd2 vssd2 vccd2 vccd2 _4211_/X sky130_fd_sc_hd__a22o_1
X_5191_ _5191_/A _5191_/B vssd2 vssd2 vccd2 vccd2 _5192_/B sky130_fd_sc_hd__xnor2_2
X_4142_ _4312_/A _4457_/B _4458_/C vssd2 vssd2 vccd2 vccd2 _4142_/X sky130_fd_sc_hd__or3_1
X_4073_ _7765_/Q _4519_/B _4519_/C vssd2 vssd2 vccd2 vccd2 _4073_/X sky130_fd_sc_hd__and3_1
XFILLER_0_92_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_13_wb_clk_i clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7804_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_7832_ _7838_/CLK _7832_/D _7591_/Y vssd2 vssd2 vccd2 vccd2 _7832_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6568__A1 _6939_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4933__A _5011_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_93_518 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4975_ _4904_/A _4904_/B _4902_/Y vssd2 vssd2 vccd2 vccd2 _4977_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_46_401 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7763_ _7800_/CLK _7763_/D _7522_/Y vssd2 vssd2 vccd2 vccd2 _7763_/Q sky130_fd_sc_hd__dfrtp_4
X_6714_ _6714_/A _6714_/B vssd2 vssd2 vccd2 vccd2 _6718_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_272 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3926_ _4252_/D _4707_/A vssd2 vssd2 vccd2 vccd2 _4030_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_46_445 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7694_ _7806_/CLK _7694_/D vssd2 vssd2 vccd2 vccd2 _7694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_520 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6645_ _6645_/A _6645_/B vssd2 vssd2 vccd2 vccd2 _6647_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_73_275 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_6_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3857_ _3888_/B _7795_/Q _7796_/Q _3860_/B vssd2 vssd2 vccd2 vccd2 _3858_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_104_517 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6576_ _6576_/A _6576_/B _6576_/C vssd2 vssd2 vccd2 vccd2 _6578_/A sky130_fd_sc_hd__or3_1
XANTENNA__6740__A1 _6668_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_26_180 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5527_ _5528_/C _5528_/D _5030_/C _4814_/Y vssd2 vssd2 vccd2 vccd2 _5529_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_41_161 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5458_ _5458_/A _5528_/B _5458_/C vssd2 vssd2 vccd2 vccd2 _5528_/C sky130_fd_sc_hd__or3_2
Xfanout200 _4257_/Y vssd2 vssd2 vccd2 vccd2 _4711_/A sky130_fd_sc_hd__buf_4
X_4409_ _4409_/A _4409_/B vssd2 vssd2 vccd2 vccd2 _4412_/A sky130_fd_sc_hd__xnor2_2
X_5389_ _5328_/A _5431_/B _5388_/X vssd2 vssd2 vccd2 vccd2 _5390_/B sky130_fd_sc_hd__o21a_2
Xfanout222 _5414_/A vssd2 vssd2 vccd2 vccd2 _5315_/B sky130_fd_sc_hd__clkbuf_8
X_7128_ _7031_/B _7031_/C _7211_/B vssd2 vssd2 vccd2 vccd2 _7128_/X sky130_fd_sc_hd__a21o_1
Xfanout255 _6253_/A vssd2 vssd2 vccd2 vccd2 _6670_/A sky130_fd_sc_hd__clkbuf_8
Xfanout233 _6358_/B vssd2 vssd2 vccd2 vccd2 _6587_/B sky130_fd_sc_hd__clkbuf_8
Xfanout244 _3913_/Y vssd2 vssd2 vccd2 vccd2 _4814_/B sky130_fd_sc_hd__buf_4
X_7059_ _7060_/A _7060_/B vssd2 vssd2 vccd2 vccd2 _7114_/A sky130_fd_sc_hd__nor2_1
Xfanout288 _7629_/A vssd2 vssd2 vccd2 vccd2 _7645_/A sky130_fd_sc_hd__buf_4
Xfanout277 _7453_/Y vssd2 vssd2 vccd2 vccd2 _7454_/C sky130_fd_sc_hd__buf_6
Xfanout266 _7806_/Q vssd2 vssd2 vccd2 vccd2 _3888_/B sky130_fd_sc_hd__buf_4
XFILLER_0_96_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4282__A2 _4044_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5939__A _7844_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_96_345 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1213 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_96_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1257 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4562__B _5276_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1268 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_592 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_52_404 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7365__S _7383_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_103_561 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6655__D _7140_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_99_161 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_62_25 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_87_378 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4760_ _4760_/A _4760_/B vssd2 vssd2 vccd2 vccd2 _4761_/B sky130_fd_sc_hd__nand2_1
X_4691_ _4691_/A _4691_/B vssd2 vssd2 vccd2 vccd2 _4693_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_43_426 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_53 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6430_ _6668_/A _6430_/B vssd2 vssd2 vccd2 vccd2 _6438_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_234 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_97 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6361_ _6357_/X _6359_/X _6281_/B vssd2 vssd2 vccd2 vccd2 _7224_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_51_470 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5312_ _5313_/B _5313_/A vssd2 vssd2 vccd2 vccd2 _5370_/A sky130_fd_sc_hd__and2b_1
X_6292_ _6294_/A _6294_/B vssd2 vssd2 vccd2 vccd2 _6292_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_87_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5243_ _5243_/A _5243_/B vssd2 vssd2 vccd2 vccd2 _5248_/A sky130_fd_sc_hd__xnor2_1
X_5174_ _5175_/B _5175_/A vssd2 vssd2 vccd2 vccd2 _5174_/Y sky130_fd_sc_hd__nand2b_1
Xhold19 hold19/A vssd2 vssd2 vccd2 vccd2 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_4125_ _7767_/Q _4125_/B _4125_/C vssd2 vssd2 vccd2 vccd2 _4125_/X sky130_fd_sc_hd__and3_1
XANTENNA__6789__A1 _6150_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4366__C _4711_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_78_312 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4056_ _7727_/D _4093_/A vssd2 vssd2 vccd2 vccd2 _4094_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_36_92 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7815_ _7826_/CLK _7815_/D _7574_/Y vssd2 vssd2 vccd2 vccd2 _7815_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_507 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_93_337 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_78_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_19_423 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4958_ _4958_/A _4958_/B vssd2 vssd2 vccd2 vccd2 _4960_/B sky130_fd_sc_hd__xor2_1
X_7746_ _7771_/CLK _7746_/D _7505_/Y vssd2 vssd2 vccd2 vccd2 _7746_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_562 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4889_ _4889_/A _4889_/B vssd2 vssd2 vccd2 vccd2 _4890_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_46_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3909_ _7787_/Q _7788_/Q vssd2 vssd2 vccd2 vccd2 _3910_/D sky130_fd_sc_hd__or2_1
X_7677_ _7806_/CLK _7677_/D vssd2 vssd2 vccd2 vccd2 _7677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_61_212 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6628_ _6670_/A _6629_/B _6629_/C vssd2 vssd2 vccd2 vccd2 _7197_/B sky130_fd_sc_hd__and3_4
XFILLER_0_6_383 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_15_673 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6559_ _6481_/A _6481_/C _6481_/B vssd2 vssd2 vccd2 vccd2 _6561_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_61_289 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_42_492 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__6475__D _7253_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_88_109 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_69_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__5452__A1 _5451_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5669__A _6283_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_96_153 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_69_378 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XTAP_1021 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_69_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1065 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5204__A1 _5404_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5204__B2 _5328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1098 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_510 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_25_426 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_108_675 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6704__A1 _6705_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_4_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6704__B2 _6783_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_40_429 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_57_25 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_805 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_849 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5930_ _6664_/A vssd2 vssd2 vccd2 vccd2 _6812_/B sky130_fd_sc_hd__inv_2
XFILLER_0_73_68 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5994__A2 _5993_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_75_326 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5861_ _6105_/A _6707_/A vssd2 vssd2 vccd2 vccd2 _5862_/B sky130_fd_sc_hd__nor2_1
X_7600_ _7627_/A vssd2 vssd2 vccd2 vccd2 _7600_/Y sky130_fd_sc_hd__inv_2
X_4812_ _5042_/B _5220_/A vssd2 vssd2 vccd2 vccd2 _4819_/A sky130_fd_sc_hd__nor2_2
X_5792_ _7845_/Q _6253_/B _6191_/C _6191_/D vssd2 vssd2 vccd2 vccd2 _5798_/B sky130_fd_sc_hd__and4_1
XFILLER_0_90_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4743_ _4656_/A _4809_/B _3827_/Y _4809_/A vssd2 vssd2 vccd2 vccd2 _4745_/B sky130_fd_sc_hd__a22o_1
X_7531_ _7564_/A vssd2 vssd2 vccd2 vccd2 _7531_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_22_61 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_71_532 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7462_ _7702_/Q _7454_/C _7485_/B1 hold253/X vssd2 vssd2 vccd2 vccd2 _7462_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3827__A _4809_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_113_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6413_ _6783_/A _7037_/A _6345_/B _6343_/Y vssd2 vssd2 vccd2 vccd2 _6422_/A sky130_fd_sc_hd__o31ai_4
XFILLER_0_71_565 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_71_554 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4674_ _4606_/A _4606_/B _4604_/X vssd2 vssd2 vccd2 vccd2 _4676_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_98_65 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7393_ _7436_/A _7393_/B vssd2 vssd2 vccd2 vccd2 _7665_/D sky130_fd_sc_hd__and2_1
XFILLER_0_24_481 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_101_317 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6344_ _6344_/A _6344_/B vssd2 vssd2 vccd2 vccd2 _6345_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_12_643 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6275_ _6812_/A _6812_/B _6989_/A _7047_/A vssd2 vssd2 vccd2 vccd2 _6276_/C sky130_fd_sc_hd__or4b_1
XANTENNA__7034__A _7034_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_51_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5226_ _5227_/A _5227_/B _5227_/C vssd2 vssd2 vccd2 vccd2 _5272_/A sky130_fd_sc_hd__a21o_1
XANTENNA__5131__B1 _5548_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5157_ _5158_/A _5158_/B vssd2 vssd2 vccd2 vccd2 _5159_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_91 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5088_ _5089_/A _5089_/B vssd2 vssd2 vccd2 vccd2 _5162_/B sky130_fd_sc_hd__nand2_1
X_4108_ _4809_/A _4082_/B _4082_/D _3995_/X _3880_/D vssd2 vssd2 vccd2 vccd2 _4108_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_78_120 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4039_ _7765_/Q _4125_/B _4125_/C _7761_/Q _4815_/B vssd2 vssd2 vccd2 vccd2 _4039_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_79_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_78_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_66_337 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_115 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_104 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_109_417 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_148 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_137 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_126 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_93_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XPHY_159 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7729_ _7793_/CLK _7729_/D _7488_/Y vssd2 vssd2 vccd2 vccd2 _7729_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_275 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_104_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5374__D _5528_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_104_177 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6783__A _6783_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_57_326 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XPHY_6 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_57_348 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_57_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_53_521 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold308 hold308/A vssd2 vssd2 vccd2 vccd2 la_data_out[31] sky130_fd_sc_hd__buf_12
XFILLER_0_53_587 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_40_226 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_111_637 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4390_ _4388_/X _4390_/B vssd2 vssd2 vccd2 vccd2 _4391_/B sky130_fd_sc_hd__nand2b_1
Xhold319 _7757_/Q vssd2 vssd2 vccd2 vccd2 hold319/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5361__B1 _5528_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_40_248 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_68_79 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XTAP_602 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _6122_/B vssd2 vssd2 vccd2 vccd2 _6184_/A sky130_fd_sc_hd__inv_2
XTAP_635 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _5011_/A _5550_/A vssd2 vssd2 vccd2 vccd2 _5012_/B sky130_fd_sc_hd__or2_1
XTAP_679 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_41 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_108_85 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_23_7 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6962_ _6897_/A _6897_/B _6895_/X vssd2 vssd2 vccd2 vccd2 _6963_/B sky130_fd_sc_hd__a21o_1
X_5913_ _5913_/A _5913_/B vssd2 vssd2 vccd2 vccd2 _5915_/B sky130_fd_sc_hd__xor2_2
X_6893_ _6893_/A _6893_/B vssd2 vssd2 vccd2 vccd2 _6896_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_48_315 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__3978__A1 _7765_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5844_ _6402_/A _5907_/D vssd2 vssd2 vccd2 vccd2 _5862_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_412 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_75_178 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_75_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_99_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_91_649 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4660__B _5468_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_44_521 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7514_ _7564_/A vssd2 vssd2 vccd2 vccd2 _7514_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_201 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5775_ _5772_/X _5774_/X _5938_/C vssd2 vssd2 vccd2 vccd2 _5775_/Y sky130_fd_sc_hd__o21ai_1
X_4726_ wire212/X _4881_/A2 _4880_/B vssd2 vssd2 vccd2 vccd2 _4728_/B sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout222_A _5414_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_16_234 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7445_ hold158/X _7803_/D _7451_/S vssd2 vssd2 vccd2 vccd2 _7445_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_640 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4657_ _4268_/A _5458_/A _4454_/B vssd2 vssd2 vccd2 vccd2 _4657_/X sky130_fd_sc_hd__o21a_1
Xinput91 input91/A vssd2 vssd2 vccd2 vccd2 input91/X sky130_fd_sc_hd__clkbuf_1
Xinput80 wbs_adr_i[8] vssd2 vssd2 vccd2 vccd2 _7341_/B sky130_fd_sc_hd__buf_1
X_7376_ _7452_/A _7376_/B vssd2 vssd2 vccd2 vccd2 _7658_/D sky130_fd_sc_hd__and2_1
XFILLER_0_102_648 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_101_125 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6327_ _6707_/A _6479_/C vssd2 vssd2 vccd2 vccd2 _6330_/C sky130_fd_sc_hd__nor2_1
X_4588_ _4585_/X _4586_/X _4519_/B vssd2 vssd2 vccd2 vccd2 _5081_/C sky130_fd_sc_hd__o21ai_4
XFILLER_0_101_169 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6258_ _6259_/A _6259_/B vssd2 vssd2 vccd2 vccd2 _6335_/A sky130_fd_sc_hd__nor2_2
X_6189_ _6189_/A _6189_/B _6188_/A vssd2 vssd2 vccd2 vccd2 _6316_/A sky130_fd_sc_hd__or3b_1
XANTENNA__6852__B1 _7222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5209_ _5210_/B _5528_/A _5498_/D _5210_/A vssd2 vssd2 vccd2 vccd2 _5211_/A sky130_fd_sc_hd__o22ai_2
XANTENNA__5781__A_N _6670_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_79_462 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_94_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_66_101 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4630__A2 _5142_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_13_19 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_109_225 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_54_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_35_510 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_62_340 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_35_565 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_50_524 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_62_395 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_50_546 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7373__S _7383_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_22_248 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6497__B _6572_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_38_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7096__B1 _7294_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_89_237 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6018__A _6670_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_281 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_85_454 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_85_443 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_85_421 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_73_605 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_70_47 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_57_156 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3890_ _7791_/Q _4162_/A _4141_/D _4100_/B vssd2 vssd2 vccd2 vccd2 _3890_/X sky130_fd_sc_hd__and4_1
XFILLER_0_45_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5560_ _5516_/A _5543_/A _5543_/B vssd2 vssd2 vccd2 vccd2 _5560_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_26_554 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4385__B2 _4809_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4511_ wire212/X _4881_/A2 _5222_/A vssd2 vssd2 vccd2 vccd2 _4513_/B sky130_fd_sc_hd__a21oi_2
X_5491_ _5456_/A _5455_/B _5455_/A vssd2 vssd2 vccd2 vccd2 _5492_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_53 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_79_78 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7230_ _7259_/B _7230_/B vssd2 vssd2 vccd2 vccd2 _7232_/C sky130_fd_sc_hd__nand2_1
X_4442_ _4402_/A _4402_/B _4400_/X vssd2 vssd2 vccd2 vccd2 _4452_/A sky130_fd_sc_hd__a21bo_2
Xhold105 _7486_/X vssd2 vssd2 vccd2 vccd2 _7726_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 wbs_adr_i[0] vssd2 vssd2 vccd2 vccd2 input50/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 input84/X vssd2 vssd2 vccd2 vccd2 hold127/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 wbs_dat_i[7] vssd2 vssd2 vccd2 vccd2 input96/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _7451_/X vssd2 vssd2 vccd2 vccd2 _7452_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_97 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7161_ _7162_/A _7162_/B vssd2 vssd2 vccd2 vccd2 _7205_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_1_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_21_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4373_ _4268_/A _4125_/B _4067_/X vssd2 vssd2 vccd2 vccd2 _4373_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_95_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6112_ _6111_/B _6111_/C _6111_/A vssd2 vssd2 vccd2 vccd2 _6112_/X sky130_fd_sc_hd__a21o_1
X_7092_ _7140_/A _7237_/A _7138_/C _7253_/B vssd2 vssd2 vccd2 vccd2 _7093_/B sky130_fd_sc_hd__or4_1
XTAP_410 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _5907_/D _5994_/X _6150_/B _6590_/A vssd2 vssd2 vccd2 vccd2 _6045_/B sky130_fd_sc_hd__a22o_1
XANTENNA__5098__C1 _4267_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_443 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7312__A _7326_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_487 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_82 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4860__A2 _5404_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_fanout172_A _6150_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1609 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_70 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6945_ _6986_/A _7181_/A vssd2 vssd2 vccd2 vccd2 _6946_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5767__A _6550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_91_413 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_76_465 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7011__B1 _6939_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_48_178 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6876_ _6876_/A _6876_/B vssd2 vssd2 vccd2 vccd2 _6885_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5827_ _6282_/A _6018_/D _5811_/B _7846_/Q _6191_/D vssd2 vssd2 vccd2 vccd2 _5827_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_91_457 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_17_554 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5758_ _6152_/B _5944_/B _7846_/Q vssd2 vssd2 vccd2 vccd2 _5759_/C sky130_fd_sc_hd__and3b_1
XANTENNA__4376__A1 _4328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4376__B2 _7770_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4709_ _4709_/A _4709_/B vssd2 vssd2 vccd2 vccd2 _4718_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__7314__A1 _7253_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7314__B2 _7253_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5689_ _5690_/B _5690_/C _7882_/Q vssd2 vssd2 vccd2 vccd2 _5691_/A sky130_fd_sc_hd__o21ai_4
X_7428_ _7436_/A _7428_/B vssd2 vssd2 vccd2 vccd2 _7682_/D sky130_fd_sc_hd__and2_1
XANTENNA__4128__A1 _7768_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5876__A1 _7843_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_32_568 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold661 hold661/A vssd2 vssd2 vccd2 vccd2 hold661/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold650 _7821_/Q vssd2 vssd2 vccd2 vccd2 hold650/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5876__B2 _7844_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_12_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xhold672 wbs_adr_i[22] vssd2 vssd2 vccd2 vccd2 input64/A sky130_fd_sc_hd__dlygate4sd3_1
X_7359_ hold207/X _7762_/D _7383_/S vssd2 vssd2 vccd2 vccd2 _7359_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_292 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold694 _7690_/Q vssd2 vssd2 vccd2 vccd2 hold694/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 _7680_/Q vssd2 vssd2 vccd2 vccd2 hold683/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7222__A _7222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_99_557 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7250__B1 _7336_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_67_410 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_24_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_79_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_67_443 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_94_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6356__A2 _5816_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_638 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_82_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_23_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_373 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_112_209 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_105_261 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_50_387 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__6816__B1 _6668_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4991_ _4920_/A _4920_/B _4918_/Y vssd2 vssd2 vccd2 vccd2 _4993_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_81_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6730_ _7037_/A _7045_/A vssd2 vssd2 vccd2 vccd2 _6731_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_58_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_58_454 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_18_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3942_ _4068_/B _3982_/B vssd2 vssd2 vccd2 vccd2 _4427_/A sky130_fd_sc_hd__nor2_4
X_6661_ _6661_/A _6661_/B vssd2 vssd2 vccd2 vccd2 _6681_/A sky130_fd_sc_hd__xor2_2
X_3873_ _3813_/A _3813_/B _4745_/A _4454_/B _4656_/C vssd2 vssd2 vccd2 vccd2 _4326_/D
+ sky130_fd_sc_hd__a2111oi_4
X_6592_ _6592_/A _6592_/B vssd2 vssd2 vccd2 vccd2 _6595_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_148 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_26_340 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5612_ _7865_/Q _5612_/B vssd2 vssd2 vccd2 vccd2 _5620_/B sky130_fd_sc_hd__xnor2_2
X_5543_ _5543_/A _5543_/B vssd2 vssd2 vccd2 vccd2 _5561_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_26_351 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_26_362 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_41_332 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5474_ _5407_/A _5407_/B _5405_/B vssd2 vssd2 vccd2 vccd2 _5476_/B sky130_fd_sc_hd__a21bo_1
X_7213_ _6767_/A _6767_/B _6767_/C _7025_/X _7211_/X vssd2 vssd2 vccd2 vccd2 _7216_/B
+ sky130_fd_sc_hd__a311o_1
X_4425_ _4405_/A _4405_/B _4403_/Y vssd2 vssd2 vccd2 vccd2 _4440_/A sky130_fd_sc_hd__a21oi_4
X_7144_ _7144_/A _7144_/B vssd2 vssd2 vccd2 vccd2 _7146_/A sky130_fd_sc_hd__nor2_1
X_4356_ _4356_/A _4356_/B vssd2 vssd2 vccd2 vccd2 _4418_/B sky130_fd_sc_hd__xnor2_2
XTAP_240 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7075_ _7075_/A _7075_/B vssd2 vssd2 vccd2 vccd2 _7077_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__4666__A _4896_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4287_ _4287_/A _4287_/B vssd2 vssd2 vccd2 vccd2 _4289_/B sky130_fd_sc_hd__xnor2_2
XTAP_262 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ _6026_/A _6026_/B vssd2 vssd2 vccd2 vccd2 _6055_/A sky130_fd_sc_hd__xor2_1
XANTENNA__7480__B1 _7483_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_295 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6586__A2 _5816_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_76_262 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6928_ _6928_/A _6928_/B vssd2 vssd2 vccd2 vccd2 _6930_/B sky130_fd_sc_hd__xor2_1
XANTENNA__6338__A2 _6571_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6859_ _6860_/A _6860_/B vssd2 vssd2 vccd2 vccd2 _6859_/X sky130_fd_sc_hd__and2_1
XFILLER_0_36_104 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_37_627 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_107_537 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_64_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_107_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_44_192 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_44_170 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_253 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5849__B2 _7844_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5849__A1 _7842_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_32_398 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_3_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold480 la_data_in[13] vssd2 vssd2 vccd2 vccd2 hold43/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 hold28/X vssd2 vssd2 vccd2 vccd2 _7886_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6274__A1 _6664_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6274__B2 _5931_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7471__B1 _7483_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_67_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6329__A2 _6404_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5001__A2 _4996_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_70_416 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_113_529 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_51_663 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_11_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_11_538 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_11_527 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_2_248 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4210_ _4328_/A _4125_/B _3931_/Y _4252_/D _7767_/Q vssd2 vssd2 vccd2 vccd2 _4210_/X
+ sky130_fd_sc_hd__a32o_1
X_5190_ _5191_/A _5191_/B vssd2 vssd2 vccd2 vccd2 _5190_/Y sky130_fd_sc_hd__nand2_1
X_4141_ _4521_/A _4458_/C _4141_/C _4141_/D vssd2 vssd2 vccd2 vccd2 _4141_/X sky130_fd_sc_hd__or4_1
XANTENNA__7462__B1 _7485_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4072_ _4058_/X _4059_/X _4065_/X _4071_/X _3965_/A vssd2 vssd2 vccd2 vccd2 _4072_/Y
+ sky130_fd_sc_hd__o41ai_2
X_7831_ _7838_/CLK _7831_/D _7590_/Y vssd2 vssd2 vccd2 vccd2 _7831_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6568__A2 _6572_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4933__B _5076_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4028__B1 _7767_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_58_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4974_ _4974_/A _4974_/B vssd2 vssd2 vccd2 vccd2 _4977_/A sky130_fd_sc_hd__xnor2_4
X_7762_ _7800_/CLK _7762_/D _7521_/Y vssd2 vssd2 vccd2 vccd2 _7762_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_86_571 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6713_ _6939_/A _7181_/A vssd2 vssd2 vccd2 vccd2 _6714_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_46_413 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_3925_ _7788_/Q _3925_/B vssd2 vssd2 vccd2 vccd2 _4063_/B sky130_fd_sc_hd__xnor2_4
X_7693_ _7804_/CLK _7693_/D vssd2 vssd2 vccd2 vccd2 _7693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_295 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6644_ _6554_/X _6558_/B _6555_/X vssd2 vssd2 vccd2 vccd2 _6645_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_46_457 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3856_ _7795_/Q _3822_/A _7796_/Q _3888_/B vssd2 vssd2 vccd2 vccd2 _3858_/A sky130_fd_sc_hd__o211ai_2
XFILLER_0_81_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6575_ _6652_/B _6574_/C _6574_/A vssd2 vssd2 vccd2 vccd2 _6576_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__6740__A2 _7313_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_61_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7037__A _7037_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5526_ _5526_/A _5528_/D vssd2 vssd2 vccd2 vccd2 _5530_/A sky130_fd_sc_hd__nor2_1
X_5457_ _5414_/B _5498_/D _4814_/Y _5326_/A vssd2 vssd2 vccd2 vccd2 _5459_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_41_184 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_112_595 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4408_ _4408_/A _4408_/B vssd2 vssd2 vccd2 vccd2 _4409_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__5780__A _6281_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout223 _4460_/X vssd2 vssd2 vccd2 vccd2 _5222_/A sky130_fd_sc_hd__clkbuf_8
X_5388_ _5388_/A _5388_/B vssd2 vssd2 vccd2 vccd2 _5388_/X sky130_fd_sc_hd__xor2_1
Xfanout201 _4257_/Y vssd2 vssd2 vccd2 vccd2 _5210_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7127_ _7023_/A _7080_/Y _7082_/B vssd2 vssd2 vccd2 vccd2 _7127_/X sky130_fd_sc_hd__a21o_1
Xfanout256 _7854_/Q vssd2 vssd2 vccd2 vccd2 _6253_/A sky130_fd_sc_hd__clkbuf_8
X_4339_ _4882_/A _4966_/A _4283_/A _4284_/Y vssd2 vssd2 vccd2 vccd2 _4348_/A sky130_fd_sc_hd__o31ai_4
X_7058_ _7058_/A _7058_/B vssd2 vssd2 vccd2 vccd2 _7060_/B sky130_fd_sc_hd__xnor2_1
Xfanout267 _4049_/B vssd2 vssd2 vccd2 vccd2 _4050_/B sky130_fd_sc_hd__buf_6
Xfanout278 _7440_/A vssd2 vssd2 vccd2 vccd2 _7436_/A sky130_fd_sc_hd__clkbuf_4
Xfanout289 _7629_/A vssd2 vssd2 vccd2 vccd2 _7627_/A sky130_fd_sc_hd__buf_8
X_6009_ _6059_/A _6064_/A vssd2 vssd2 vccd2 vccd2 _6010_/B sky130_fd_sc_hd__nand2_1
XTAP_1214 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_357 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1247 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_287 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_52_416 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_17_192 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_103_573 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__6786__A _7047_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7381__S _7383_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_16_608 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_83_574 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_55_265 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4690_ _4551_/A _4551_/B _4619_/C _4688_/X _4689_/X vssd2 vssd2 vccd2 vccd2 _4691_/B
+ sky130_fd_sc_hd__o311a_4
XFILLER_0_43_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_36_490 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_113_337 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_102_65 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_11_52 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6360_ _6357_/X _6359_/X _6281_/B vssd2 vssd2 vccd2 vccd2 _7099_/B sky130_fd_sc_hd__o21a_4
XFILLER_0_51_482 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_11_302 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5311_ _5276_/A _5528_/A _5550_/B _5210_/B vssd2 vssd2 vccd2 vccd2 _5313_/B sky130_fd_sc_hd__o22a_1
X_6291_ _6668_/A _7047_/A _6229_/B _6227_/X vssd2 vssd2 vccd2 vccd2 _6294_/B sky130_fd_sc_hd__a31o_1
X_5242_ _5242_/A _5242_/B vssd2 vssd2 vccd2 vccd2 _5243_/B sky130_fd_sc_hd__xor2_2
X_5173_ _5175_/A _5175_/B vssd2 vssd2 vccd2 vccd2 _5173_/X sky130_fd_sc_hd__and2b_1
X_4124_ _4162_/A _4251_/B vssd2 vssd2 vccd2 vccd2 _4124_/X sky130_fd_sc_hd__and2_1
XANTENNA__6789__A2 _7145_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4366__D _4782_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xinput1 input1/A vssd2 vssd2 vccd2 vccd2 input1/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4249__B1 _7766_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4055_ _4898_/A _4882_/A vssd2 vssd2 vccd2 vccd2 _4093_/A sky130_fd_sc_hd__or2_1
XFILLER_0_78_324 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_93_305 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7814_ _7814_/CLK _7814_/D _7573_/Y vssd2 vssd2 vccd2 vccd2 _7814_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_109 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_93_349 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4957_ _4958_/A _4958_/B vssd2 vssd2 vccd2 vccd2 _5024_/A sky130_fd_sc_hd__and2b_1
X_7745_ _7771_/CLK _7745_/D _7504_/Y vssd2 vssd2 vccd2 vccd2 _7745_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_435 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_19_457 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_74_585 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4888_ _4889_/A _4889_/B vssd2 vssd2 vccd2 vccd2 _4949_/B sky130_fd_sc_hd__and2_1
X_7676_ _7806_/CLK _7676_/D vssd2 vssd2 vccd2 vccd2 _7676_/Q sky130_fd_sc_hd__dfxtp_1
X_3908_ _7783_/Q _7784_/Q _7785_/Q _7786_/Q vssd2 vssd2 vccd2 vccd2 _3910_/C sky130_fd_sc_hd__or4_2
XFILLER_0_19_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6627_ _6627_/A _6627_/B vssd2 vssd2 vccd2 vccd2 _6627_/X sky130_fd_sc_hd__xor2_1
X_3839_ _3813_/A _3813_/B _4458_/D _4144_/C _4326_/C vssd2 vssd2 vccd2 vccd2 _4267_/C
+ sky130_fd_sc_hd__a2111oi_2
XANTENNA__4724__A1 _4810_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6558_ _6558_/A _6558_/B vssd2 vssd2 vccd2 vccd2 _6561_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_373 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6489_ _6489_/A _6489_/B vssd2 vssd2 vccd2 vccd2 _6491_/B sky130_fd_sc_hd__xnor2_2
X_5509_ _5510_/A _5510_/B vssd2 vssd2 vccd2 vccd2 _5541_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_100_521 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_10_390 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5988__B1 _7845_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_96_121 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5452__A2 _5451_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1022 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_165 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1044 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5204__A2 _5414_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_32_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XTAP_1099 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4963__B2 _4962_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_92_382 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_80_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_65_596 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_52_235 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_52_224 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_577 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6704__A2 _7253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_52_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_460 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_40_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_110_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_817 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_549 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7405__A _7452_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_839 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7140__A _7140_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6275__D_N _7047_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5860_ _5857_/X _5858_/X _5859_/X _5734_/Y vssd2 vssd2 vccd2 vccd2 _5860_/Y sky130_fd_sc_hd__o31ai_1
X_4811_ _4811_/A _4811_/B vssd2 vssd2 vccd2 vccd2 _4822_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_56_541 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5791_ _6253_/B _6253_/C _6191_/D vssd2 vssd2 vccd2 vccd2 _5791_/X sky130_fd_sc_hd__and3_1
X_4742_ _4742_/A _4803_/A vssd2 vssd2 vccd2 vccd2 _4748_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_585 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_56_563 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7530_ _7565_/A vssd2 vssd2 vccd2 vccd2 _7530_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_276 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4673_ _4673_/A _4673_/B vssd2 vssd2 vccd2 vccd2 _4676_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_511 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_43_202 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7461_ _7701_/Q _7454_/C _7485_/B1 hold235/X vssd2 vssd2 vccd2 vccd2 _7461_/X sky130_fd_sc_hd__a22o_1
X_6412_ _6412_/A _6412_/B vssd2 vssd2 vccd2 vccd2 _6450_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__6203__B _7037_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_43_257 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_98_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_71_599 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_71_588 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_43_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7392_ hold187/X _7665_/Q _7418_/S vssd2 vssd2 vccd2 vccd2 _7392_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4706__B2 _4809_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_24_460 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4004__A _4454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_113_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_101_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6343_ _6344_/A _6344_/B vssd2 vssd2 vccd2 vccd2 _6343_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_51_290 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6274_ _6664_/A _6150_/B _6571_/C _5931_/C vssd2 vssd2 vccd2 vccd2 _6276_/B sky130_fd_sc_hd__a22o_1
X_5225_ _5225_/A _5225_/B vssd2 vssd2 vccd2 vccd2 _5227_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__5131__A1 _5133_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_44_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5156_ _5156_/A _5156_/B vssd2 vssd2 vccd2 vccd2 _5158_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_70 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6873__B _7253_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5087_ _5087_/A _5087_/B vssd2 vssd2 vccd2 vccd2 _5089_/B sky130_fd_sc_hd__xor2_1
X_4107_ _4105_/X _4106_/X _3993_/D vssd2 vssd2 vccd2 vccd2 _4115_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_611 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7050__A _7143_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4038_ _3987_/X _4028_/X _4037_/X _4033_/C _4035_/X vssd2 vssd2 vccd2 vccd2 _4044_/A
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_78_154 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_93_113 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_66_305 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_116 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_109_429 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_94_658 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XPHY_149 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_138 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_66_349 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_127 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_47_541 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5989_ _6158_/A _5937_/B _5935_/D _6283_/A vssd2 vssd2 vccd2 vccd2 _5989_/X sky130_fd_sc_hd__a22o_1
X_7728_ _7776_/CLK _7728_/D _7487_/Y vssd2 vssd2 vccd2 vccd2 _7728_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_254 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_62_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7659_ _7787_/CLK _7659_/D vssd2 vssd2 vccd2 vccd2 _7659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_408 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_34_246 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_62_599 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_15_482 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_15_493 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_30_441 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_104_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_100_351 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_30_496 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4881__B1 _5498_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6783__B _7255_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_441 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4633__B1 _4782_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_485 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XPHY_7 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_72_319 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_65_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_53_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_38_596 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_108_495 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_80_385 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_80_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_25_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold309 hold662/X vssd2 vssd2 vccd2 vccd2 hold663/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5361__B2 _5404_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5361__A1 _5081_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_111_649 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_68_36 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_603 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5008_/X _5010_/B vssd2 vssd2 vccd2 vccd2 _5012_/A sky130_fd_sc_hd__and2b_1
XTAP_636 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_53 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4494__A _4898_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_17_40 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_17_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_108_97 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6961_ _6961_/A _6961_/B vssd2 vssd2 vccd2 vccd2 _6963_/A sky130_fd_sc_hd__xnor2_2
X_5912_ _5913_/A _5913_/B vssd2 vssd2 vccd2 vccd2 _5962_/A sky130_fd_sc_hd__nand2_1
X_6892_ _6891_/B _6891_/C _6891_/A vssd2 vssd2 vccd2 vccd2 _6893_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_113 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5843_ _6550_/A _6092_/A vssd2 vssd2 vccd2 vccd2 _5863_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_33_50 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_91_617 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_29_552 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_29_574 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_33_72 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7513_ _7641_/A vssd2 vssd2 vccd2 vccd2 _7513_/Y sky130_fd_sc_hd__inv_2
X_5774_ _7845_/Q _5937_/B _5935_/D _7847_/Q vssd2 vssd2 vccd2 vccd2 _5774_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_71_352 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4725_ _5029_/A _5315_/B vssd2 vssd2 vccd2 vccd2 _4728_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_114_421 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7444_ _7452_/A _7444_/B vssd2 vssd2 vccd2 vccd2 _7444_/X sky130_fd_sc_hd__and2_1
X_4656_ _4656_/A _4656_/B _4656_/C vssd2 vssd2 vccd2 vccd2 _4656_/X sky130_fd_sc_hd__or3_1
XFILLER_0_12_430 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7375_ hold107/X _7658_/Q _7383_/S vssd2 vssd2 vccd2 vccd2 _7375_/X sky130_fd_sc_hd__mux2_1
Xinput81 wbs_adr_i[9] vssd2 vssd2 vccd2 vccd2 _7341_/A sky130_fd_sc_hd__clkbuf_1
Xinput70 wbs_adr_i[28] vssd2 vssd2 vccd2 vccd2 input70/X sky130_fd_sc_hd__clkbuf_1
X_4587_ _4585_/X _4586_/X _4519_/B vssd2 vssd2 vccd2 vccd2 _5326_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_101_137 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6326_ _6550_/A _7181_/A vssd2 vssd2 vccd2 vccd2 _6332_/A sky130_fd_sc_hd__nor2_1
XANTENNA__7045__A _7045_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_12_452 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xinput92 input92/A vssd2 vssd2 vccd2 vccd2 input92/X sky130_fd_sc_hd__clkbuf_1
X_6257_ _6550_/A _7051_/A vssd2 vssd2 vccd2 vccd2 _6259_/B sky130_fd_sc_hd__or2_1
X_6188_ _6188_/A _6188_/B vssd2 vssd2 vccd2 vccd2 _7815_/D sky130_fd_sc_hd__xnor2_1
X_5208_ _5208_/A _5208_/B vssd2 vssd2 vccd2 vccd2 _5217_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__6852__A1 _6039_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5139_ _5139_/A _5139_/B vssd2 vssd2 vccd2 vccd2 _5139_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_8_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7723_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_603 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4091__A1 _4598_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_39_305 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_94_444 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_349 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_109_237 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_94_499 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_47_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_35_500 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_62_352 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_50_558 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_15_290 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7096__A1 _7143_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_30_260 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7096__B2 _7143_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_38_39 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_89_205 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_89_249 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_58_603 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_57_102 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_97_293 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_85_433 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_70_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_26_511 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_26_522 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_38_360 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_38_371 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_53_341 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5873__A _7845_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_26_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4510_ _5029_/A _5099_/A vssd2 vssd2 vccd2 vccd2 _4513_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_53_374 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5490_ _5490_/A _5490_/B vssd2 vssd2 vccd2 vccd2 _5492_/A sky130_fd_sc_hd__or2_1
XFILLER_0_102_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4441_ _4441_/A _4441_/B vssd2 vssd2 vccd2 vccd2 _4471_/A sky130_fd_sc_hd__xor2_4
Xhold117 _7351_/X vssd2 vssd2 vccd2 vccd2 _7420_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold106 wbs_dat_i[11] vssd2 vssd2 vccd2 vccd2 input85/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_558 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_110_65 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7160_ _7045_/A _7255_/B _7095_/A _7093_/B vssd2 vssd2 vccd2 vccd2 _7162_/B sky130_fd_sc_hd__o31a_1
Xhold128 _7408_/X vssd2 vssd2 vccd2 vccd2 _7409_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_644 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold139 input96/X vssd2 vssd2 vccd2 vccd2 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
X_6111_ _6111_/A _6111_/B _6111_/C vssd2 vssd2 vccd2 vccd2 _6111_/Y sky130_fd_sc_hd__nand3_1
X_4372_ _4372_/A _4372_/B vssd2 vssd2 vccd2 vccd2 _4409_/A sky130_fd_sc_hd__xnor2_2
XTAP_400 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_271 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7091_ _6430_/B _7222_/A _7222_/C _7197_/A vssd2 vssd2 vccd2 vccd2 _7093_/A sky130_fd_sc_hd__a22o_1
XTAP_411 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_293 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6042_ _6039_/X _6040_/X _5992_/B vssd2 vssd2 vccd2 vccd2 _6989_/A sky130_fd_sc_hd__o21ai_4
XTAP_444 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6944_ _6944_/A _6944_/B vssd2 vssd2 vccd2 vccd2 _6946_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_433 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_76_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7011__B2 _7291_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6875_ _6927_/A _6875_/B vssd2 vssd2 vccd2 vccd2 _6875_/X sky130_fd_sc_hd__and2_1
X_5826_ _6158_/A _5826_/B vssd2 vssd2 vccd2 vccd2 _5826_/X sky130_fd_sc_hd__and2_1
XFILLER_0_17_500 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_91_447 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5757_ _5992_/B _5992_/C _5757_/C vssd2 vssd2 vccd2 vccd2 _5760_/C sky130_fd_sc_hd__and3b_1
XANTENNA__6879__A _6973_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4708_ _4708_/A _5550_/A vssd2 vssd2 vccd2 vccd2 _4709_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5783__A _6093_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_8_298 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__7314__A2 _7291_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5688_ _5735_/B _7881_/Q vssd2 vssd2 vccd2 vccd2 _5690_/C sky130_fd_sc_hd__and2_1
X_7427_ hold207/X _7794_/D _7451_/S vssd2 vssd2 vccd2 vccd2 _7427_/X sky130_fd_sc_hd__mux2_1
X_4639_ _4639_/A _4639_/B vssd2 vssd2 vccd2 vccd2 _4640_/B sky130_fd_sc_hd__xnor2_1
Xhold640 _7834_/Q vssd2 vssd2 vccd2 vccd2 hold640/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 _7831_/Q vssd2 vssd2 vccd2 vccd2 hold662/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 hold651/A vssd2 vssd2 vccd2 vccd2 hold651/X sky130_fd_sc_hd__dlygate4sd3_1
X_7358_ _7436_/A _7358_/B vssd2 vssd2 vccd2 vccd2 _7649_/D sky130_fd_sc_hd__and2_1
X_6309_ _6387_/A _6320_/B vssd2 vssd2 vccd2 vccd2 _6310_/B sky130_fd_sc_hd__or2_1
X_7289_ _7289_/A _7289_/B vssd2 vssd2 vccd2 vccd2 _7290_/B sky130_fd_sc_hd__or2_1
Xhold673 _7340_/X vssd2 vssd2 vccd2 vccd2 _7346_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 _7662_/Q vssd2 vssd2 vccd2 vccd2 hold695/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 _7688_/Q vssd2 vssd2 vccd2 vccd2 hold684/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7222__B _7222_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_219 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4064__A1 _7763_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4064__B2 _7765_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_39_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__5013__B1 _5081_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_54_149 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_23_514 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_2_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_23_536 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_23_558 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4846__A_N _4769_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_35_385 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_105_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_50_399 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_49_38 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6816__B2 _6669_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7413__A _7452_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3941__A _7767_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4990_ _4990_/A _4990_/B vssd2 vssd2 vccd2 vccd2 _4993_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_58_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_14_52 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3941_ _7767_/Q _4814_/B _4315_/B _4214_/B vssd2 vssd2 vccd2 vccd2 _3941_/X sky130_fd_sc_hd__and4_1
X_6660_ _6660_/A _6660_/B vssd2 vssd2 vccd2 vccd2 _6661_/B sky130_fd_sc_hd__xnor2_2
X_3872_ _3813_/A _3813_/B _4454_/B vssd2 vssd2 vccd2 vccd2 _4002_/A sky130_fd_sc_hd__a21oi_2
X_6591_ _6591_/A _6591_/B vssd2 vssd2 vccd2 vccd2 _6592_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_609 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_45_138 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5611_ _7865_/Q _5612_/B vssd2 vssd2 vccd2 vccd2 _6191_/D sky130_fd_sc_hd__xor2_4
X_5542_ _5541_/A _5541_/B _5541_/C vssd2 vssd2 vccd2 vccd2 _5543_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_480 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_5_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_30_51 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5473_ _5473_/A _5473_/B vssd2 vssd2 vccd2 vccd2 _5478_/A sky130_fd_sc_hd__nor2_1
X_7212_ _7029_/A _7029_/B _7211_/X vssd2 vssd2 vccd2 vccd2 _7216_/A sky130_fd_sc_hd__a21o_1
X_4424_ _4424_/A _4424_/B vssd2 vssd2 vccd2 vccd2 _7735_/D sky130_fd_sc_hd__xor2_1
X_7143_ _7143_/A _7143_/B _7294_/C _7313_/B vssd2 vssd2 vccd2 vccd2 _7144_/B sky130_fd_sc_hd__and4_1
X_4355_ _4355_/A _4355_/B vssd2 vssd2 vccd2 vccd2 _4356_/B sky130_fd_sc_hd__xor2_2
X_7074_ _7075_/A _7075_/B vssd2 vssd2 vccd2 vccd2 _7125_/A sky130_fd_sc_hd__nor2_1
XTAP_230 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4666__B _5220_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4286_ _4287_/B _4287_/A vssd2 vssd2 vccd2 vccd2 _4323_/A sky130_fd_sc_hd__and2b_1
XTAP_263 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _6026_/A _6026_/B vssd2 vssd2 vccd2 vccd2 _6119_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5491__B1 _5455_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_296 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout282_A _7563_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XTAP_1429 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_580 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_49_422 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6927_ _6927_/A _6927_/B vssd2 vssd2 vccd2 vccd2 _6928_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_49_488 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_9_541 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6858_ _6221_/X _6223_/X _6152_/B _7143_/A vssd2 vssd2 vccd2 vccd2 _6860_/B sky130_fd_sc_hd__o211a_1
XFILLER_0_107_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__6105__C _6989_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_9_574 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5809_ _7850_/Q _5812_/C _5920_/D _5807_/X vssd2 vssd2 vccd2 vccd2 _5809_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_36_138 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6402__A _6402_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6789_ _6150_/B _7145_/A _6785_/X _6787_/Y vssd2 vssd2 vccd2 vccd2 _6790_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_51_108 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_32_355 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_221 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_102_265 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold470 input47/X vssd2 vssd2 vccd2 vccd2 hold8/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 hold43/X vssd2 vssd2 vccd2 vccd2 input5/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 la_data_in[42] vssd2 vssd2 vccd2 vccd2 hold61/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4576__B _5099_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6274__A2 _6150_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_208 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7379__S _7383_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4037__A1 _4162_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_95_561 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_51_17 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_55_403 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_82_222 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_82_266 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_63_491 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_23_311 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_50_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_11_517 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__7143__A _7143_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4140_ _4807_/A _4863_/A vssd2 vssd2 vccd2 vccd2 _4229_/A sky130_fd_sc_hd__nor2_1
X_4071_ _4454_/A _4029_/X _4066_/X _4069_/X _4070_/X vssd2 vssd2 vccd2 vccd2 _4071_/X
+ sky130_fd_sc_hd__a2111o_1
X_7830_ _7838_/CLK _7830_/D _7589_/Y vssd2 vssd2 vccd2 vccd2 _7830_/Q sky130_fd_sc_hd__dfrtp_1
X_4973_ _4973_/A _4973_/B vssd2 vssd2 vccd2 vccd2 _4974_/B sky130_fd_sc_hd__xor2_4
X_7761_ _7795_/CLK _7761_/D _7520_/Y vssd2 vssd2 vccd2 vccd2 _7761_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5776__A1 _7843_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6712_ _6712_/A _6712_/B vssd2 vssd2 vccd2 vccd2 _6714_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_46_425 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_18_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3924_ _7788_/Q _3925_/B vssd2 vssd2 vccd2 vccd2 _4707_/A sky130_fd_sc_hd__xor2_4
X_7692_ _7804_/CLK _7692_/D vssd2 vssd2 vccd2 vccd2 _7692_/Q sky130_fd_sc_hd__dfxtp_1
X_6643_ _6643_/A _6643_/B vssd2 vssd2 vccd2 vccd2 _6645_/A sky130_fd_sc_hd__xnor2_1
X_3855_ _7793_/Q _7792_/Q _7791_/Q _7794_/Q _3888_/B vssd2 vssd2 vccd2 vccd2 _3860_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_0_33_108 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6574_ _6574_/A _6652_/B _6574_/C vssd2 vssd2 vccd2 vccd2 _6576_/B sky130_fd_sc_hd__and3_1
XFILLER_0_61_439 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7037__B _7253_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5525_ _5525_/A _5525_/B vssd2 vssd2 vccd2 vccd2 _7753_/D sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_22_wb_clk_i clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7739_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5456_ _5456_/A _5456_/B vssd2 vssd2 vccd2 vccd2 _7751_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_563 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4407_ _4407_/A _4407_/B vssd2 vssd2 vccd2 vccd2 _4408_/B sky130_fd_sc_hd__xor2_4
XANTENNA__7053__A _7237_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5387_ _5388_/A _5388_/B vssd2 vssd2 vccd2 vccd2 _5439_/A sky130_fd_sc_hd__and2b_1
Xfanout213 _6404_/D vssd2 vssd2 vccd2 vccd2 _7143_/B sky130_fd_sc_hd__clkbuf_8
Xfanout202 _4217_/Y vssd2 vssd2 vccd2 vccd2 _4662_/B sky130_fd_sc_hd__buf_4
X_7126_ _7126_/A _7126_/B vssd2 vssd2 vccd2 vccd2 _7211_/C sky130_fd_sc_hd__nand2_2
X_4338_ _4338_/A _4338_/B vssd2 vssd2 vccd2 vccd2 _4350_/A sky130_fd_sc_hd__xnor2_4
Xfanout246 _3830_/X vssd2 vssd2 vccd2 vccd2 _4458_/D sky130_fd_sc_hd__clkbuf_8
Xfanout224 _4460_/X vssd2 vssd2 vccd2 vccd2 _5431_/A sky130_fd_sc_hd__buf_2
Xfanout235 _6191_/C vssd2 vssd2 vccd2 vccd2 _6253_/C sky130_fd_sc_hd__clkbuf_4
X_7057_ _7057_/A _7057_/B vssd2 vssd2 vccd2 vccd2 _7058_/B sky130_fd_sc_hd__xor2_1
X_4269_ _4809_/A _4268_/D _4002_/B _7766_/Q _4656_/C vssd2 vssd2 vccd2 vccd2 _4269_/X
+ sky130_fd_sc_hd__a32o_1
Xfanout279 _7450_/A vssd2 vssd2 vccd2 vccd2 _7440_/A sky130_fd_sc_hd__clkbuf_4
Xfanout268 _7774_/Q vssd2 vssd2 vccd2 vccd2 _4809_/A sky130_fd_sc_hd__buf_6
Xfanout257 _7853_/Q vssd2 vssd2 vccd2 vccd2 _6510_/A sky130_fd_sc_hd__buf_4
X_6008_ _6008_/A _6008_/B vssd2 vssd2 vccd2 vccd2 _6064_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_69_528 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XTAP_1204 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1248 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_241 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1259 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_583 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_64_211 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_92_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_64_244 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__5519__A1 _5451_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_107_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_60_450 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_32_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__6786__B _7094_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_68_583 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_55_233 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_28_436 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__7138__A _7237_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_70_214 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_55_288 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_3_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_113_305 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_102_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_113_349 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6290_ _6290_/A _6290_/B vssd2 vssd2 vccd2 vccd2 _6294_/A sky130_fd_sc_hd__xnor2_2
X_5310_ _5357_/C _5310_/B vssd2 vssd2 vccd2 vccd2 _7748_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_163 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7132__B1 _7034_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_51_494 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5241_ _5187_/A _5187_/B _5185_/Y vssd2 vssd2 vccd2 vccd2 _5242_/B sky130_fd_sc_hd__a21o_1
X_5172_ _5101_/A _5101_/B _5099_/X vssd2 vssd2 vccd2 vccd2 _5175_/B sky130_fd_sc_hd__a21bo_1
X_4123_ _4328_/A _4057_/X _4121_/X _3971_/Y _4122_/X vssd2 vssd2 vccd2 vccd2 _4123_/X
+ sky130_fd_sc_hd__a221o_1
Xinput2 input2/A vssd2 vssd2 vccd2 vccd2 input2/X sky130_fd_sc_hd__clkbuf_1
X_4054_ _5455_/A _4096_/A vssd2 vssd2 vccd2 vccd2 _4095_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4249__A1 _4893_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7601__A _7627_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_36_72 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7813_ _7814_/CLK _7813_/D _7572_/Y vssd2 vssd2 vccd2 vccd2 _7813_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_317 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7744_ _7771_/CLK _7744_/D _7503_/Y vssd2 vssd2 vccd2 vccd2 _7744_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_594 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4956_ _4956_/A _4956_/B vssd2 vssd2 vccd2 vccd2 _4958_/B sky130_fd_sc_hd__xor2_1
X_4887_ _4887_/A _4887_/B vssd2 vssd2 vccd2 vccd2 _4889_/B sky130_fd_sc_hd__xor2_1
X_7675_ _7787_/CLK _7675_/D vssd2 vssd2 vccd2 vccd2 _7675_/Q sky130_fd_sc_hd__dfxtp_1
X_3907_ _7783_/Q _7784_/Q vssd2 vssd2 vccd2 vccd2 _3907_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_406 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6626_ _6626_/A vssd2 vssd2 vccd2 vccd2 _6758_/A sky130_fd_sc_hd__inv_2
XFILLER_0_74_597 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_6_330 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3838_ _7799_/Q _3838_/B vssd2 vssd2 vccd2 vccd2 _4144_/D sky130_fd_sc_hd__xnor2_2
XANTENNA__4724__A2 _4880_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6557_ _6783_/A _7181_/A vssd2 vssd2 vccd2 vccd2 _6558_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_42_461 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_14_152 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5508_ _5478_/A _5478_/B _5473_/A vssd2 vssd2 vccd2 vccd2 _5510_/B sky130_fd_sc_hd__a21oi_1
X_6488_ _6488_/A _6488_/B vssd2 vssd2 vccd2 vccd2 _6489_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_30_645 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_100_533 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5439_ _5439_/A _5439_/B vssd2 vssd2 vccd2 vccd2 _5440_/B sky130_fd_sc_hd__or2_1
XANTENNA__4488__A1 _7771_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4200__A _4268_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4488__B2 _7772_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7109_ _7109_/A _7109_/B vssd2 vssd2 vccd2 vccd2 _7111_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__7511__A _7564_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5988__A1 _6253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5669__C _6424_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_96_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XTAP_1012 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_96_177 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1045 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4963__A2 _5406_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_37_244 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_37_266 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_80_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_52_247 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7392__S _7418_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3923__B1 _4050_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_33_483 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XTAP_807 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4110__A _7767_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_88_601 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_87_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_73_48 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7140__B _7255_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4810_ _4810_/A _5498_/D vssd2 vssd2 vccd2 vccd2 _4811_/B sky130_fd_sc_hd__or2_2
XFILLER_0_68_391 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_56_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_8_628 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5790_ _6157_/A _6071_/B _6019_/C _5921_/D vssd2 vssd2 vccd2 vccd2 _5798_/A sky130_fd_sc_hd__and4_1
XTAP_1590 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_83_361 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4741_ _4962_/A _5164_/A _4965_/B _5406_/A vssd2 vssd2 vccd2 vccd2 _4803_/A sky130_fd_sc_hd__or4_1
XFILLER_0_56_575 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4672_ _4672_/A _4672_/B vssd2 vssd2 vccd2 vccd2 _4673_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_56_597 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7460_ _7700_/Q _7454_/C _7485_/B1 hold239/X vssd2 vssd2 vccd2 vccd2 _7460_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_22_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_114_625 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_113_113 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6411_ _6411_/A _6411_/B vssd2 vssd2 vccd2 vccd2 _6412_/B sky130_fd_sc_hd__xor2_4
XANTENNA__5903__A1 _6282_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_31_409 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7391_ _7436_/A _7391_/B vssd2 vssd2 vccd2 vccd2 _7664_/D sky130_fd_sc_hd__and2_1
XANTENNA__5903__B2 _6157_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_24_472 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6342_ _6939_/A _6973_/A vssd2 vssd2 vccd2 vccd2 _6344_/B sky130_fd_sc_hd__nor2_2
X_6273_ _6581_/A _6939_/A vssd2 vssd2 vccd2 vccd2 _6276_/A sky130_fd_sc_hd__nor2_1
X_5224_ _5224_/A _5224_/B vssd2 vssd2 vccd2 vccd2 _5225_/B sky130_fd_sc_hd__xnor2_1
X_5155_ _5082_/A _5084_/B _5082_/B vssd2 vssd2 vccd2 vccd2 _5156_/B sky130_fd_sc_hd__a21boi_2
XANTENNA_fanout195_A _5207_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5086_ _5087_/A _5087_/B vssd2 vssd2 vccd2 vccd2 _5162_/A sky130_fd_sc_hd__nand2_1
X_4106_ _7763_/Q _4809_/B _4146_/B _7764_/Q vssd2 vssd2 vccd2 vccd2 _4106_/X sky130_fd_sc_hd__a22o_1
XANTENNA__7050__B _7222_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4037_ _4162_/A _4427_/A _4164_/C _4036_/X _4021_/X vssd2 vssd2 vccd2 vccd2 _4037_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_94_637 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_78_188 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_106 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_93_125 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_128 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_117 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5988_ _6253_/A _5850_/B _5936_/B _7845_/Q _6510_/B vssd2 vssd2 vccd2 vccd2 _5988_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_93_169 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4939_ _5210_/B _5222_/A _5315_/B _5210_/A vssd2 vssd2 vccd2 vccd2 _4941_/A sky130_fd_sc_hd__o22ai_1
X_7727_ _7776_/CLK _7727_/D _7436_/A vssd2 vssd2 vccd2 vccd2 _7727_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_244 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_62_523 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7658_ _7787_/CLK _7658_/D vssd2 vssd2 vccd2 vccd2 _7658_/Q sky130_fd_sc_hd__dfxtp_1
X_6609_ _6610_/A _6610_/B _6610_/C vssd2 vssd2 vccd2 vccd2 _6694_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_62_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_6_160 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7589_ _7590_/A vssd2 vssd2 vccd2 vccd2 _7589_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4849__B _4849_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_30_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_100_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_97_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4633__A1 _4711_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4633__B2 _4966_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_85_615 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_69_177 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_69_155 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_8 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_72_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_93_670 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_25_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4105__A _7766_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_108_485 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_53_556 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_53_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_40_206 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5361__A2 _5498_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_68_59 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_21_497 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_604 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4494__B _5276_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_108_65 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6960_ _6960_/A _6960_/B vssd2 vssd2 vccd2 vccd2 _6961_/B sky130_fd_sc_hd__nor2_1
X_5911_ _6402_/A _5907_/D _5862_/B _5863_/B _5863_/A vssd2 vssd2 vccd2 vccd2 _5913_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_8 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_76_626 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_48_306 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6891_ _6891_/A _6891_/B _6891_/C vssd2 vssd2 vccd2 vccd2 _6893_/A sky130_fd_sc_hd__and3_1
XFILLER_0_75_125 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5842_ _5826_/X _5832_/X _5838_/X _5840_/X _5665_/B vssd2 vssd2 vccd2 vccd2 _6092_/A
+ sky130_fd_sc_hd__o41ai_4
XFILLER_0_75_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_63_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4388__B1 _5042_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_8_436 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5773_ _6152_/B _5944_/B _6155_/B vssd2 vssd2 vccd2 vccd2 _5935_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_33_84 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_90_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_84_670 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4724_ _4810_/A _4880_/B _4664_/B _4663_/B vssd2 vssd2 vccd2 vccd2 _4732_/A sky130_fd_sc_hd__o31a_1
X_7512_ _7564_/A vssd2 vssd2 vccd2 vccd2 _7512_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_447 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_114_433 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4655_ _4655_/A _4655_/B vssd2 vssd2 vccd2 vccd2 _4673_/A sky130_fd_sc_hd__xnor2_1
X_7443_ hold107/X _7690_/Q _7451_/S vssd2 vssd2 vccd2 vccd2 _7443_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_477 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7374_ _7452_/A _7374_/B vssd2 vssd2 vccd2 vccd2 _7657_/D sky130_fd_sc_hd__and2_1
Xinput82 wbs_cyc_i vssd2 vssd2 vccd2 vccd2 _7453_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput71 wbs_adr_i[29] vssd2 vssd2 vccd2 vccd2 input71/X sky130_fd_sc_hd__clkbuf_1
Xinput60 wbs_adr_i[19] vssd2 vssd2 vccd2 vccd2 _7344_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_291 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_31_228 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4586_ _4809_/A _4519_/C _4146_/B _4268_/A vssd2 vssd2 vccd2 vccd2 _4586_/X sky130_fd_sc_hd__a22o_1
XANTENNA_fanout208_A _4704_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_101_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__7045__B _7140_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_12_442 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xinput93 input93/A vssd2 vssd2 vccd2 vccd2 input93/X sky130_fd_sc_hd__buf_1
X_6325_ _6071_/X _6323_/X _6016_/B vssd2 vssd2 vccd2 vccd2 _6642_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_101_149 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_12_497 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6256_ _7143_/B vssd2 vssd2 vccd2 vccd2 _7051_/A sky130_fd_sc_hd__inv_2
XFILLER_0_58_81 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6187_ _6189_/A _6189_/B _6069_/A vssd2 vssd2 vccd2 vccd2 _6188_/B sky130_fd_sc_hd__o21a_1
X_5207_ _5207_/A _5550_/A vssd2 vssd2 vccd2 vccd2 _5208_/B sky130_fd_sc_hd__nor2_1
XANTENNA__6852__A2 _6040_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5138_ _5139_/A _5139_/B vssd2 vssd2 vccd2 vccd2 _5243_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_442 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5069_ _5069_/A _5133_/C vssd2 vssd2 vccd2 vccd2 _7744_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__4091__A2 _4807_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_66_125 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_66_114 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_109_205 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_54_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_109_249 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_81_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_556 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7096__A2 _7222_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_38_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_89_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_97_261 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_57_136 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6359__B2 _6093_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6359__A1 _6253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_70_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5031__A1 _5030_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_38_383 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_72_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_53_353 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_183 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_53_386 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4440_ _4440_/A _4440_/B vssd2 vssd2 vccd2 vccd2 _4441_/B sky130_fd_sc_hd__xnor2_4
Xhold107 input85/X vssd2 vssd2 vccd2 vccd2 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
Xhold129 _7409_/X vssd2 vssd2 vccd2 vccd2 _7673_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 _7352_/X vssd2 vssd2 vccd2 vccd2 _7383_/S sky130_fd_sc_hd__buf_6
X_6110_ _6109_/A _6109_/B _6109_/C vssd2 vssd2 vccd2 vccd2 _6111_/C sky130_fd_sc_hd__a21o_1
XANTENNA__6985__A _7047_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4371_ _4372_/B _4372_/A vssd2 vssd2 vccd2 vccd2 _4475_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_95_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7090_ _7058_/A _7058_/B _7056_/X vssd2 vssd2 vccd2 vccd2 _7107_/A sky130_fd_sc_hd__a21o_1
XTAP_412 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6039_/X _6040_/X _5992_/B vssd2 vssd2 vccd2 vccd2 _6150_/B sky130_fd_sc_hd__o21a_4
XTAP_434 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_50 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6943_ _6944_/A _6944_/B vssd2 vssd2 vccd2 vccd2 _6943_/Y sky130_fd_sc_hd__nand2_1
X_6874_ _6738_/A _7294_/C _6872_/X vssd2 vssd2 vccd2 vccd2 _6875_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_44_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_48_158 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5825_ _6253_/C _6075_/C _6075_/D vssd2 vssd2 vccd2 vccd2 _5825_/X sky130_fd_sc_hd__and3_1
XFILLER_0_29_383 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_8_288 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5756_ _6158_/A _5781_/B _5850_/D _6283_/A vssd2 vssd2 vccd2 vccd2 _5757_/C sky130_fd_sc_hd__a22o_1
XANTENNA__6879__B _6973_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4781__B1 _4965_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5687_ _7881_/Q _5690_/B vssd2 vssd2 vccd2 vccd2 _5937_/B sky130_fd_sc_hd__xor2_4
X_4707_ _4707_/A _4707_/B vssd2 vssd2 vccd2 vccd2 _5145_/B sky130_fd_sc_hd__nand2_2
X_4638_ _4639_/B _4639_/A vssd2 vssd2 vccd2 vccd2 _4638_/X sky130_fd_sc_hd__and2b_1
X_7426_ _7436_/A _7426_/B vssd2 vssd2 vccd2 vccd2 _7681_/D sky130_fd_sc_hd__and2_1
Xhold630 _7816_/Q vssd2 vssd2 vccd2 vccd2 hold630/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold641 hold641/A vssd2 vssd2 vccd2 vccd2 hold641/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 hold663/A vssd2 vssd2 vccd2 vccd2 hold663/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 _7823_/Q vssd2 vssd2 vccd2 vccd2 hold652/X sky130_fd_sc_hd__dlygate4sd3_1
X_4569_ _4569_/A _4569_/B vssd2 vssd2 vccd2 vccd2 _4570_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_12_272 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7357_ hold187/X _7761_/D _7383_/S vssd2 vssd2 vccd2 vccd2 _7357_/X sky130_fd_sc_hd__mux2_1
X_6308_ _6308_/A _6308_/B vssd2 vssd2 vccd2 vccd2 _6320_/B sky130_fd_sc_hd__nor2_1
X_7288_ _7289_/A _7289_/B vssd2 vssd2 vccd2 vccd2 _7319_/A sky130_fd_sc_hd__nand2_1
Xhold696 _7689_/Q vssd2 vssd2 vccd2 vccd2 hold696/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 _7686_/Q vssd2 vssd2 vccd2 vccd2 hold685/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 _7346_/Y vssd2 vssd2 vccd2 vccd2 hold674/X sky130_fd_sc_hd__dlygate4sd3_1
X_6239_ _6173_/A _6173_/B _6171_/Y vssd2 vssd2 vccd2 vccd2 _6241_/B sky130_fd_sc_hd__o21a_1
XANTENNA__7222__C _7222_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_990 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6135__A _6572_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5261__A1 _5145_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_39_103 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_94_253 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_67_467 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_82_437 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5013__A1 _5210_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5013__B2 _4711_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_90_481 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_62_172 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_23_526 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_31_581 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_81_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_3940_ _7782_/Q _3940_/B vssd2 vssd2 vccd2 vccd2 _4214_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_105_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_58_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_18_309 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_3871_ _4656_/B _5458_/A vssd2 vssd2 vccd2 vccd2 _4103_/B sky130_fd_sc_hd__nand2_2
XANTENNA__5884__A _6158_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6590_ _6590_/A _6591_/A _7313_/B vssd2 vssd2 vccd2 vccd2 _6590_/X sky130_fd_sc_hd__and3_1
X_5610_ _5586_/B _5584_/Y _5587_/X _5599_/B vssd2 vssd2 vccd2 vccd2 _6191_/C sky130_fd_sc_hd__o211a_1
XFILLER_0_109_580 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_5_236 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_5_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_14_504 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5541_ _5541_/A _5541_/B _5541_/C vssd2 vssd2 vccd2 vccd2 _5543_/A sky130_fd_sc_hd__or3_1
XFILLER_0_26_397 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_30_63 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7211_ _7211_/A _7211_/B _7211_/C _7211_/D vssd2 vssd2 vccd2 vccd2 _7211_/X sky130_fd_sc_hd__or4_1
XFILLER_0_53_194 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_30_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5472_ _5472_/A _5472_/B _5472_/C vssd2 vssd2 vccd2 vccd2 _5473_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_41_356 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4423_ _4309_/B _4362_/B _5455_/A vssd2 vssd2 vccd2 vccd2 _4424_/B sky130_fd_sc_hd__o21a_1
X_7142_ _7143_/B _7294_/C _7313_/B _7143_/A vssd2 vssd2 vccd2 vccd2 _7144_/A sky130_fd_sc_hd__a22oi_2
XANTENNA__7604__A _7627_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_1_464 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4354_ _4355_/A _4355_/B vssd2 vssd2 vccd2 vccd2 _4354_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_39_50 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7073_ _7012_/B _7012_/C _7012_/A vssd2 vssd2 vccd2 vccd2 _7075_/B sky130_fd_sc_hd__o21ba_1
XTAP_231 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_61 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6024_ _6550_/A _6973_/A vssd2 vssd2 vccd2 vccd2 _6026_/B sky130_fd_sc_hd__nor2_1
X_4285_ _4285_/A _4285_/B vssd2 vssd2 vccd2 vccd2 _4287_/B sky130_fd_sc_hd__xor2_2
XTAP_264 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7480__A2 _7483_/A2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_297 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_529 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_68_209 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1419 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_434 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6926_ _6927_/A _6927_/B vssd2 vssd2 vccd2 vccd2 _6926_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_76_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_76_220 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_71_81 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6857_ _6152_/X _6153_/X _6159_/X _7143_/B _5944_/B vssd2 vssd2 vccd2 vccd2 _6860_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_91_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6788_ _6989_/A _6788_/B _7181_/A _6785_/X vssd2 vssd2 vccd2 vccd2 _6790_/A sky130_fd_sc_hd__or4b_1
X_5808_ _5586_/B _5584_/Y _5586_/Y _5811_/C vssd2 vssd2 vccd2 vccd2 _5920_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_9_564 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5739_ _5739_/A _5755_/C _5762_/B vssd2 vssd2 vccd2 vccd2 _5739_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__6402__B _7145_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_17_397 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4203__A _4328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_102_233 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7409_ _7452_/A _7409_/B vssd2 vssd2 vccd2 vccd2 _7409_/X sky130_fd_sc_hd__and2_1
XFILLER_0_32_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_277 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7514__A _7564_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold460 la_data_in[9] vssd2 vssd2 vccd2 vccd2 hold35/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 hold8/X vssd2 vssd2 vccd2 vccd2 _7879_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 hold61/X vssd2 vssd2 vccd2 vccd2 input37/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 input5/X vssd2 vssd2 vccd2 vccd2 hold44/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7471__A2 _7483_/A2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6431__B1 _7224_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_95_573 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_27_106 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_55_437 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_139 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_82_289 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_35_183 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_50_120 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_51_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_76_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7424__A _7436_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_76_48 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7143__B _7143_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7462__A2 _7454_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4070_ _4328_/A _4315_/B _4214_/B _4070_/D vssd2 vssd2 vccd2 vccd2 _4070_/X sky130_fd_sc_hd__and4_1
XANTENNA__5879__A _6282_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_25_63 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4972_ _4973_/A _4973_/B vssd2 vssd2 vccd2 vccd2 _4972_/Y sky130_fd_sc_hd__nor2_1
X_7760_ _7795_/CLK _7760_/D _7519_/Y vssd2 vssd2 vccd2 vccd2 _7760_/Q sky130_fd_sc_hd__dfrtp_1
X_6711_ _6989_/A _7051_/A _6712_/B vssd2 vssd2 vccd2 vccd2 _6711_/X sky130_fd_sc_hd__or3_1
XFILLER_0_58_253 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7691_ _7787_/CLK _7691_/D vssd2 vssd2 vccd2 vccd2 _7691_/Q sky130_fd_sc_hd__dfxtp_1
X_3923_ _7787_/Q _3954_/C _3910_/B _3910_/C _4050_/B vssd2 vssd2 vccd2 vccd2 _3925_/B
+ sky130_fd_sc_hd__o41a_4
X_6642_ _6855_/A _6642_/B vssd2 vssd2 vccd2 vccd2 _6643_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_18_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3854_ _7794_/Q _3854_/B vssd2 vssd2 vccd2 vccd2 _4103_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_673 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6573_ _6572_/C _6572_/D _6150_/B _6657_/B vssd2 vssd2 vccd2 vccd2 _6574_/C sky130_fd_sc_hd__a2bb2o_1
X_5524_ _5456_/A _5455_/B _5492_/A hold404/X vssd2 vssd2 vccd2 vccd2 _5525_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_14_356 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_112_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5455_ _5455_/A _5455_/B vssd2 vssd2 vccd2 vccd2 _5456_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_153 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_67_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_4406_ _4407_/A _4407_/B vssd2 vssd2 vccd2 vccd2 _4470_/A sky130_fd_sc_hd__nand2_2
X_7125_ _7125_/A _7125_/B _7125_/C vssd2 vssd2 vccd2 vccd2 _7126_/B sky130_fd_sc_hd__or3_1
XANTENNA__7053__B _7181_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout203 _4217_/Y vssd2 vssd2 vccd2 vccd2 _5164_/A sky130_fd_sc_hd__clkbuf_4
Xfanout214 _6404_/C vssd2 vssd2 vccd2 vccd2 _7143_/A sky130_fd_sc_hd__clkbuf_8
X_5386_ _5316_/A _5318_/B _5316_/B vssd2 vssd2 vccd2 vccd2 _5388_/B sky130_fd_sc_hd__a21bo_1
Xfanout225 _6549_/Y vssd2 vssd2 vccd2 vccd2 _7255_/B sky130_fd_sc_hd__clkbuf_8
X_4337_ _4337_/A _4337_/B vssd2 vssd2 vccd2 vccd2 _4338_/B sky130_fd_sc_hd__nand2_2
Xfanout236 _5588_/Y vssd2 vssd2 vccd2 vccd2 _7313_/A sky130_fd_sc_hd__buf_4
X_7056_ _7057_/A _7057_/B vssd2 vssd2 vccd2 vccd2 _7056_/X sky130_fd_sc_hd__and2_1
Xfanout258 _7853_/Q vssd2 vssd2 vccd2 vccd2 _6398_/A sky130_fd_sc_hd__clkbuf_4
X_4268_ _4268_/A _4326_/B _4326_/C _4268_/D vssd2 vssd2 vccd2 vccd2 _4268_/X sky130_fd_sc_hd__and4_1
Xfanout269 hold407/X vssd2 vssd2 vccd2 vccd2 _4893_/A sky130_fd_sc_hd__buf_8
X_6007_ _6005_/X _6007_/B vssd2 vssd2 vccd2 vccd2 _6008_/B sky130_fd_sc_hd__and2b_1
XANTENNA__4693__A _4693_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4199_ _4656_/A _3995_/X _4075_/B _4162_/A _4198_/X vssd2 vssd2 vccd2 vccd2 _4199_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_1205 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_80 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1216 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _6909_/A _6909_/B vssd2 vssd2 vccd2 vccd2 _7033_/C sky130_fd_sc_hd__and2_1
XTAP_1249 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_521 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_9_361 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5519__A2 _5451_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_24_109 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_92_598 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5029__A _5029_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4868__A _5042_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_60_462 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_32_175 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_33_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6786__C _7143_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold290 hold290/A vssd2 vssd2 vccd2 vccd2 la_data_out[27] sky130_fd_sc_hd__buf_12
XFILLER_0_46_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_87_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_68_551 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_68_573 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_83_532 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5140__A1_N _5011_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7419__A _7452_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_256 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_55_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__7138__B _7224_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_113_317 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_51_462 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5240_ _5240_/A _5240_/B vssd2 vssd2 vccd2 vccd2 _5242_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_11_348 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_11_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_87_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_11_359 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5171_ _5171_/A _5171_/B vssd2 vssd2 vccd2 vccd2 _5175_/A sky130_fd_sc_hd__xnor2_1
X_4122_ _4454_/A _4214_/C _4125_/C _4122_/D vssd2 vssd2 vccd2 vccd2 _4122_/X sky130_fd_sc_hd__and4_1
X_4053_ _7727_/D _4053_/B vssd2 vssd2 vccd2 vccd2 _4096_/A sky130_fd_sc_hd__or2_1
Xinput3 input3/A vssd2 vssd2 vccd2 vccd2 input3/X sky130_fd_sc_hd__clkbuf_1
X_7812_ _7814_/CLK _7812_/D _7571_/Y vssd2 vssd2 vccd2 vccd2 _7812_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4955_ _4956_/A _4956_/B vssd2 vssd2 vccd2 vccd2 _5035_/A sky130_fd_sc_hd__and2_1
X_7743_ _7771_/CLK _7743_/D _7502_/Y vssd2 vssd2 vccd2 vccd2 _7743_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_521 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_74_510 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_46_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3906_ _7779_/Q _7780_/Q _7781_/Q _7782_/Q vssd2 vssd2 vccd2 vccd2 _3910_/B sky130_fd_sc_hd__or4_4
X_4886_ _4887_/A _4887_/B vssd2 vssd2 vccd2 vccd2 _4949_/A sky130_fd_sc_hd__nor2_1
X_7674_ _7802_/CLK _7674_/D vssd2 vssd2 vccd2 vccd2 _7674_/Q sky130_fd_sc_hd__dfxtp_1
X_6625_ _6627_/A _6627_/B vssd2 vssd2 vccd2 vccd2 _6626_/A sky130_fd_sc_hd__and2_1
XFILLER_0_61_215 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3837_ _7799_/Q _3838_/B vssd2 vssd2 vccd2 vccd2 _4326_/C sky130_fd_sc_hd__xor2_4
XFILLER_0_34_418 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6556_ _6556_/A _6556_/B vssd2 vssd2 vccd2 vccd2 _6558_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_473 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5507_ _5539_/B _5507_/B vssd2 vssd2 vccd2 vccd2 _5510_/A sky130_fd_sc_hd__or2_1
XFILLER_0_100_501 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6487_ _6488_/A _6488_/B vssd2 vssd2 vccd2 vccd2 _6566_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_42_484 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_2_570 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5438_ _5439_/A _5439_/B vssd2 vssd2 vccd2 vccd2 _5486_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_100_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5369_ _5370_/A _5370_/B _5370_/C vssd2 vssd2 vccd2 vccd2 _5430_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_100_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7108_ _7109_/A _7109_/B vssd2 vssd2 vccd2 vccd2 _7158_/A sky130_fd_sc_hd__nand2_1
X_7039_ _7153_/A _7039_/B vssd2 vssd2 vccd2 vccd2 _7042_/A sky130_fd_sc_hd__and2_1
XFILLER_0_69_337 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1013 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XTAP_1035 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_510 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_107_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_80_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_37_256 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_108_645 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_92_395 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_92_362 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_25_418 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_37_278 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_18_492 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_33_440 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__5373__B1 _5528_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_110_309 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4598__A _4598_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_60_292 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_60_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_808 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5222__A _5222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4939__B1 _5315_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1591 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1580 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _5164_/A _4965_/B _5406_/A _4807_/A vssd2 vssd2 vccd2 vccd2 _4742_/A sky130_fd_sc_hd__o22ai_1
XFILLER_0_83_373 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4671_ _4672_/A _4672_/B vssd2 vssd2 vccd2 vccd2 _4671_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_524 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_43_215 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_16_418 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6410_ _6410_/A _6410_/B vssd2 vssd2 vccd2 vccd2 _6411_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__5892__A _6550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_43_237 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7390_ hold175/X _7776_/D _7418_/S vssd2 vssd2 vccd2 vccd2 _7390_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_637 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_113_125 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6341_ _6855_/A _6973_/B vssd2 vssd2 vccd2 vccd2 _6344_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_113_169 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6272_ _6272_/A _6272_/B vssd2 vssd2 vccd2 vccd2 _6299_/A sky130_fd_sc_hd__xor2_2
X_5223_ _5224_/A _5224_/B vssd2 vssd2 vccd2 vccd2 _5223_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_11_178 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_11_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7612__A _7613_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5154_ _5154_/A _5154_/B vssd2 vssd2 vccd2 vccd2 _5156_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__5131__A3 _5133_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4105_ _7766_/Q _4519_/B _4519_/C vssd2 vssd2 vccd2 vccd2 _4105_/X sky130_fd_sc_hd__and3_1
X_5085_ _5328_/A _5366_/A _5013_/X _5015_/B vssd2 vssd2 vccd2 vccd2 _5087_/B sky130_fd_sc_hd__o31ai_2
XFILLER_0_47_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5132__A _5133_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_78_101 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4036_ _4315_/B _4036_/B vssd2 vssd2 vccd2 vccd2 _4036_/X sky130_fd_sc_hd__and2_1
XFILLER_0_78_134 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_2_74 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_107 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_93_137 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_129 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_59_381 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_118 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5987_ _6157_/A _6281_/B _5700_/Y _6283_/B _7846_/Q vssd2 vssd2 vccd2 vccd2 _5987_/X
+ sky130_fd_sc_hd__a32o_1
X_4938_ _4938_/A _4938_/B vssd2 vssd2 vccd2 vccd2 _4947_/A sky130_fd_sc_hd__xnor2_1
X_7726_ _7758_/CLK _7726_/D vssd2 vssd2 vccd2 vccd2 _7726_/Q sky130_fd_sc_hd__dfxtp_1
X_4869_ _4869_/A _4869_/B vssd2 vssd2 vccd2 vccd2 _4872_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_513 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_47_576 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7657_ _7802_/CLK _7657_/D vssd2 vssd2 vccd2 vccd2 _7657_/Q sky130_fd_sc_hd__dfxtp_1
X_6608_ _6608_/A _6608_/B vssd2 vssd2 vccd2 vccd2 _6610_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_568 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_34_259 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7588_ _7590_/A vssd2 vssd2 vccd2 vccd2 _7588_/Y sky130_fd_sc_hd__inv_2
X_6539_ _6539_/A _6618_/B vssd2 vssd2 vccd2 vccd2 _7820_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_30_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_100_375 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__4330__A1 _7771_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6138__A _6138_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5042__A _5042_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_410 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4633__A2 _5042_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_123 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5830__B2 _7843_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XPHY_9 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_108_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_80_365 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5897__A1 _7843_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_7_19 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5897__B2 _7844_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_33_270 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_33_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_104_670 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_110_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_21_487 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_605 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7432__A _7436_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_627 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_108_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_88_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5910_ _5910_/A _5910_/B vssd2 vssd2 vccd2 vccd2 _5913_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_17_75 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_88_465 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6890_ _6932_/A _6888_/X _6818_/Y _6822_/A vssd2 vssd2 vccd2 vccd2 _6891_/C sky130_fd_sc_hd__o211ai_2
XFILLER_0_75_137 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5841_ _5826_/X _5832_/X _5838_/X _5840_/X _5665_/B vssd2 vssd2 vccd2 vccd2 _6150_/A
+ sky130_fd_sc_hd__o41a_2
XANTENNA__4388__B2 _4962_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4388__A1 _5042_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5772_ _5845_/B _5898_/C _5772_/C vssd2 vssd2 vccd2 vccd2 _5772_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_29_565 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4723_ _4651_/A _4651_/B _4648_/Y vssd2 vssd2 vccd2 vccd2 _4733_/A sky130_fd_sc_hd__o21ai_1
X_7511_ _7564_/A vssd2 vssd2 vccd2 vccd2 _7511_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_204 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7607__A _7613_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7442_ _7452_/A _7442_/B vssd2 vssd2 vccd2 vccd2 _7689_/D sky130_fd_sc_hd__and2_1
XFILLER_0_114_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4654_ _4654_/A _4654_/B vssd2 vssd2 vccd2 vccd2 _4655_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__5888__A1 _7843_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_44_568 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_12_410 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xinput61 hold97/X vssd2 vssd2 vccd2 vccd2 hold98/A sky130_fd_sc_hd__clkbuf_1
X_7373_ hold127/X _7769_/D _7383_/S vssd2 vssd2 vccd2 vccd2 _7373_/X sky130_fd_sc_hd__mux2_1
Xinput50 input50/A vssd2 vssd2 vccd2 vccd2 _7347_/B sky130_fd_sc_hd__clkbuf_1
Xinput72 input72/A vssd2 vssd2 vccd2 vccd2 input72/X sky130_fd_sc_hd__clkbuf_1
X_4585_ _4454_/A _4656_/C _4328_/B _4656_/A vssd2 vssd2 vccd2 vccd2 _4585_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_114_489 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7045__C _7253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xinput94 input94/A vssd2 vssd2 vccd2 vccd2 input94/X sky130_fd_sc_hd__clkbuf_1
Xinput83 input83/A vssd2 vssd2 vccd2 vccd2 input83/X sky130_fd_sc_hd__clkbuf_1
X_6324_ _6071_/X _6323_/X _6016_/B vssd2 vssd2 vccd2 vccd2 _7145_/A sky130_fd_sc_hd__o21a_4
X_6255_ _6252_/X _6253_/X _6254_/X _6191_/D vssd2 vssd2 vccd2 vccd2 _6404_/D sky130_fd_sc_hd__o31a_4
XANTENNA__4966__A _4966_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5206_ _5206_/A _5206_/B vssd2 vssd2 vccd2 vccd2 _5208_/A sky130_fd_sc_hd__nand2_1
X_6186_ _6186_/A _6186_/B vssd2 vssd2 vccd2 vccd2 _6188_/A sky130_fd_sc_hd__xnor2_1
X_5137_ _5077_/A _5079_/B _5077_/B vssd2 vssd2 vccd2 vccd2 _5139_/B sky130_fd_sc_hd__a21bo_1
X_5068_ _5068_/A _5128_/B vssd2 vssd2 vccd2 vccd2 _5133_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_79_432 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4019_ _4815_/B _4063_/B vssd2 vssd2 vccd2 vccd2 _4019_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__4076__B1 _7764_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_109_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_94_457 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_47_351 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7709_ _7787_/CLK _7709_/D vssd2 vssd2 vccd2 vccd2 _7709_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__7517__A _7564_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_62_365 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_35_568 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_62_387 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_15_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7398__S _7418_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_57_148 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5567__B1 _5550_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4116__A _4747_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_72_129 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5031__A2 _5030_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_79_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_41_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold108 _7443_/X vssd2 vssd2 vccd2 vccd2 _7444_/B sky130_fd_sc_hd__dlygate4sd3_1
X_4370_ _4370_/A _4441_/A _4370_/C vssd2 vssd2 vccd2 vccd2 _4372_/B sky130_fd_sc_hd__or3_1
Xhold119 _7375_/X vssd2 vssd2 vccd2 vccd2 _7376_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6985__B _7222_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_413 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_435 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6283_/A _5785_/X _6037_/X _6587_/B vssd2 vssd2 vccd2 vccd2 _6040_/X sky130_fd_sc_hd__a22o_4
XTAP_468 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_96 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_21_7 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_88_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6506__A _6581_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6942_ _6281_/X _6284_/X _5937_/B _7143_/A vssd2 vssd2 vccd2 vccd2 _6944_/B sky130_fd_sc_hd__o211a_1
X_6873_ _6873_/A _7253_/C _6872_/X vssd2 vssd2 vccd2 vccd2 _6927_/A sky130_fd_sc_hd__or3b_1
Xclkbuf_leaf_16_wb_clk_i clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7782_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_446 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5824_ _5824_/A _5824_/B vssd2 vssd2 vccd2 vccd2 _7808_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_91_405 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_209 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_60_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5755_ _5781_/B _5755_/B _5755_/C vssd2 vssd2 vccd2 vccd2 _5850_/D sky130_fd_sc_hd__nor3_1
XANTENNA__3865__A _7761_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6879__C _7224_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4781__B2 _5210_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4781__A1 _5210_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_71_151 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_44_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5686_ _7881_/Q _5690_/B vssd2 vssd2 vccd2 vccd2 _6155_/B sky130_fd_sc_hd__xnor2_4
X_4706_ _4706_/A1 _4815_/B _4427_/A _4809_/A vssd2 vssd2 vccd2 vccd2 _4707_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_114_253 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4637_ _4566_/A _4566_/B _4565_/B vssd2 vssd2 vccd2 vccd2 _4639_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_71_173 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7425_ hold187/X _7793_/D _7451_/S vssd2 vssd2 vccd2 vccd2 _7425_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_527 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_32_549 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xhold620 _7810_/Q vssd2 vssd2 vccd2 vccd2 hold620/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 _7833_/Q vssd2 vssd2 vccd2 vccd2 hold642/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 hold653/A vssd2 vssd2 vccd2 vccd2 hold653/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 hold631/A vssd2 vssd2 vccd2 vccd2 hold631/X sky130_fd_sc_hd__dlygate4sd3_1
X_4568_ _4569_/A _4569_/B vssd2 vssd2 vccd2 vccd2 _4568_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_69_92 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_12_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7356_ _7436_/A _7356_/B vssd2 vssd2 vccd2 vccd2 _7648_/D sky130_fd_sc_hd__and2_1
Xhold664 _7832_/Q vssd2 vssd2 vccd2 vccd2 hold664/X sky130_fd_sc_hd__dlygate4sd3_1
X_6307_ _6307_/A _6307_/B vssd2 vssd2 vccd2 vccd2 _6387_/B sky130_fd_sc_hd__xor2_2
X_4499_ _4436_/A _4433_/Y _4435_/B vssd2 vssd2 vccd2 vccd2 _4500_/B sky130_fd_sc_hd__a21o_1
X_7287_ _7256_/A _7256_/B _7254_/B vssd2 vssd2 vccd2 vccd2 _7289_/B sky130_fd_sc_hd__a21bo_1
Xhold686 _7685_/Q vssd2 vssd2 vccd2 vccd2 hold686/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 _7758_/Q vssd2 vssd2 vccd2 vccd2 hold697/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 _7789_/Q vssd2 vssd2 vccd2 vccd2 _3927_/A sky130_fd_sc_hd__buf_1
X_6238_ _6238_/A _6238_/B vssd2 vssd2 vccd2 vccd2 _6241_/A sky130_fd_sc_hd__xor2_2
XANTENNA__7483__B1 _7483_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6169_ _6169_/A _6169_/B vssd2 vssd2 vccd2 vccd2 _6172_/A sky130_fd_sc_hd__xnor2_2
XTAP_980 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_516 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_991 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7222__D _7294_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6038__A1 _7846_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6038__B2 _6253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6416__A _6939_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_79_240 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5261__A2 _5431_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_94_221 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_94_265 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_82_416 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5013__A2 _5414_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_67_479 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_54_107 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_75_490 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_35_343 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_90_493 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_90_471 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_62_162 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_62_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_50_346 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__7474__B1 _7483_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7226__B1 _6669_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6326__A _6550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5788__B1 _5736_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_81_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_45_107 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3870_ _4745_/A _4656_/C vssd2 vssd2 vccd2 vccd2 _3892_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_66_490 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5540_ _5558_/A _5540_/B vssd2 vssd2 vccd2 vccd2 _5541_/C sky130_fd_sc_hd__and2_1
XFILLER_0_26_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_53_173 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_26_387 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5471_ _5472_/A _5472_/B _5472_/C vssd2 vssd2 vccd2 vccd2 _5473_/A sky130_fd_sc_hd__o21a_1
X_7210_ _7210_/A _7210_/B vssd2 vssd2 vccd2 vccd2 _7279_/A sky130_fd_sc_hd__and2_1
X_4422_ _4422_/A _4422_/B vssd2 vssd2 vccd2 vccd2 _4424_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__6996__A _7140_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_111_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_41_368 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7141_ _7141_/A _7141_/B vssd2 vssd2 vccd2 vccd2 _7152_/A sky130_fd_sc_hd__xnor2_2
X_4353_ _4294_/A _4294_/B _4292_/X vssd2 vssd2 vccd2 vccd2 _4355_/B sky130_fd_sc_hd__a21oi_2
X_7072_ _7072_/A _7072_/B vssd2 vssd2 vccd2 vccd2 _7075_/A sky130_fd_sc_hd__xnor2_1
X_4284_ _4285_/A _4285_/B vssd2 vssd2 vccd2 vccd2 _4284_/Y sky130_fd_sc_hd__nand2b_1
XTAP_232 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7465__B1 _7485_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_254 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_95 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6023_ _6020_/X _6021_/X _5811_/B vssd2 vssd2 vccd2 vccd2 _6973_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__6105__D_N _7047_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_298 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout170_A _6138_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1409 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6925_ _6925_/A _6925_/B vssd2 vssd2 vccd2 vccd2 _6927_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_232 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_49_446 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6856_ _6856_/A _6856_/B vssd2 vssd2 vccd2 vccd2 _6866_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6787_ _7047_/A _7094_/A _7143_/A _7143_/B vssd2 vssd2 vccd2 vccd2 _6787_/Y sky130_fd_sc_hd__nand4_1
X_3999_ _7763_/Q _4328_/B vssd2 vssd2 vccd2 vccd2 _3999_/Y sky130_fd_sc_hd__nand2_1
X_5807_ _6253_/A _6194_/B _5807_/C vssd2 vssd2 vccd2 vccd2 _5807_/X sky130_fd_sc_hd__and3_1
XFILLER_0_91_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5738_ _5691_/A _5691_/B _6152_/B _5944_/B _5937_/B vssd2 vssd2 vccd2 vccd2 _6102_/C
+ sky130_fd_sc_hd__a2111oi_2
XFILLER_0_72_493 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_72_460 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_44_184 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5669_ _6283_/A _7855_/Q _6424_/A vssd2 vssd2 vccd2 vccd2 _5669_/X sky130_fd_sc_hd__and3_1
XFILLER_0_102_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7408_ hold127/X _7673_/Q _7418_/S vssd2 vssd2 vccd2 vccd2 _7408_/X sky130_fd_sc_hd__mux2_1
Xmax_cap180 _6986_/A vssd2 vssd2 vccd2 vccd2 _7045_/A sky130_fd_sc_hd__clkbuf_4
Xhold450 input30/X vssd2 vssd2 vccd2 vccd2 hold20/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 hold35/X vssd2 vssd2 vccd2 vccd2 input48/A sky130_fd_sc_hd__dlygate4sd3_1
X_7339_ _7339_/A _7339_/B _7339_/C _7339_/D vssd2 vssd2 vccd2 vccd2 _7339_/X sky130_fd_sc_hd__or4_1
Xhold472 la_data_in[18] vssd2 vssd2 vccd2 vccd2 hold41/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_289 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold494 input37/X vssd2 vssd2 vccd2 vccd2 hold62/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 hold44/X vssd2 vssd2 vccd2 vccd2 _7884_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7456__B1 _7485_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5315__A _5404_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_99_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_99_357 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6431__A1 _5816_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_95_585 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_82_213 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_106_584 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_50_132 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_31_390 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_76_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7143__C _7294_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7440__A _7440_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_92_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_25_42 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_86_541 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4433__B1 _4782_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_58_243 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_4971_ _4900_/A _4900_/B _4898_/X vssd2 vssd2 vccd2 vccd2 _4973_/B sky130_fd_sc_hd__a21boi_4
XFILLER_0_86_563 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6710_ _7047_/A _7143_/A vssd2 vssd2 vccd2 vccd2 _6712_/B sky130_fd_sc_hd__nand2_1
X_7690_ _7802_/CLK _7690_/D vssd2 vssd2 vccd2 vccd2 _7690_/Q sky130_fd_sc_hd__dfxtp_1
X_3922_ _7787_/Q _3922_/B vssd2 vssd2 vccd2 vccd2 _4253_/B sky130_fd_sc_hd__xor2_2
X_6641_ _6641_/A _6641_/B vssd2 vssd2 vccd2 vccd2 _6643_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3853_ _7794_/Q _3854_/B vssd2 vssd2 vccd2 vccd2 _3993_/D sky130_fd_sc_hd__xor2_4
XFILLER_0_27_652 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6572_ _6989_/A _6572_/B _6572_/C _6572_/D vssd2 vssd2 vccd2 vccd2 _6652_/B sky130_fd_sc_hd__or4_1
XFILLER_0_73_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_54_482 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5523_ _5544_/B _5523_/B vssd2 vssd2 vccd2 vccd2 _5525_/A sky130_fd_sc_hd__and2_1
XFILLER_0_26_184 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_41_110 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7615__A _7641_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5454_ _5454_/A _5454_/B _5547_/C vssd2 vssd2 vccd2 vccd2 _5455_/B sky130_fd_sc_hd__or3b_1
X_4405_ _4405_/A _4405_/B vssd2 vssd2 vccd2 vccd2 _4407_/B sky130_fd_sc_hd__xor2_4
X_5385_ _5385_/A _5385_/B vssd2 vssd2 vccd2 vccd2 _5390_/A sky130_fd_sc_hd__xnor2_4
X_7124_ _7125_/A _7125_/B _7125_/C vssd2 vssd2 vccd2 vccd2 _7126_/A sky130_fd_sc_hd__o21ai_2
X_4336_ _4863_/A _4662_/B _4336_/C vssd2 vssd2 vccd2 vccd2 _4337_/B sky130_fd_sc_hd__or3_1
Xfanout204 _4207_/Y vssd2 vssd2 vccd2 vccd2 _4966_/A sky130_fd_sc_hd__clkbuf_8
Xfanout237 _5164_/B vssd2 vssd2 vccd2 vccd2 _5498_/D sky130_fd_sc_hd__buf_4
Xfanout259 _7852_/Q vssd2 vssd2 vccd2 vccd2 _6093_/A sky130_fd_sc_hd__clkbuf_8
X_4267_ _4656_/A _4519_/C _4267_/C _4267_/D vssd2 vssd2 vccd2 vccd2 _4267_/X sky130_fd_sc_hd__and4_1
Xfanout248 _4809_/B vssd2 vssd2 vccd2 vccd2 _4656_/C sky130_fd_sc_hd__clkbuf_8
X_7055_ _7140_/A _7181_/A _6997_/A _6994_/Y vssd2 vssd2 vccd2 vccd2 _7057_/B sky130_fd_sc_hd__o31ai_2
X_6006_ _6003_/Y _6004_/X _5955_/Y _5960_/A vssd2 vssd2 vccd2 vccd2 _6007_/B sky130_fd_sc_hd__a211o_1
X_4198_ _4454_/A _4326_/B _4326_/C _4268_/D vssd2 vssd2 vccd2 vccd2 _4198_/X sky130_fd_sc_hd__and4_1
XANTENNA__6413__A1 _6783_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1239 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_92 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1217 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_541 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6908_ _6908_/A _6908_/B vssd2 vssd2 vccd2 vccd2 _7033_/B sky130_fd_sc_hd__xnor2_2
X_6839_ _6839_/A _6839_/B vssd2 vssd2 vccd2 vccd2 _7025_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_37_449 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_107_337 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_52_408 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_9_373 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5029__B _5498_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4868__B _5276_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_60_474 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7525__A _7557_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6786__D _7143_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold280 hold280/A vssd2 vssd2 vccd2 vccd2 la_data_out[9] sky130_fd_sc_hd__buf_12
Xhold291 hold650/X vssd2 vssd2 vccd2 vccd2 hold651/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4884__A _5030_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_305 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_95_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_83_566 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_55_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_11_33 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4124__A _4162_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_113_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_70_238 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_51_441 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_11_44 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_87_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_11_327 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5170_ _5171_/A _5171_/B vssd2 vssd2 vccd2 vccd2 _5227_/B sky130_fd_sc_hd__or2_1
X_4121_ _4122_/D _4066_/C _4120_/X _4252_/D _7765_/Q vssd2 vssd2 vccd2 vccd2 _4121_/X
+ sky130_fd_sc_hd__a32o_1
X_4052_ _4052_/A _4052_/B vssd2 vssd2 vccd2 vccd2 _7728_/D sky130_fd_sc_hd__xor2_1
XANTENNA__5402__B _5547_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xinput4 input4/A vssd2 vssd2 vccd2 vccd2 input4/X sky130_fd_sc_hd__buf_1
XFILLER_0_78_338 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7811_ _7814_/CLK _7811_/D _7570_/Y vssd2 vssd2 vccd2 vccd2 _7811_/Q sky130_fd_sc_hd__dfrtp_1
X_4954_ _5030_/A _5030_/B _4954_/C vssd2 vssd2 vccd2 vccd2 _4956_/B sky130_fd_sc_hd__and3_1
X_7742_ _7787_/CLK _7742_/D _7501_/Y vssd2 vssd2 vccd2 vccd2 _7742_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3905_ _7776_/Q _7775_/Q _7777_/Q _7778_/Q vssd2 vssd2 vccd2 vccd2 _3954_/C sky130_fd_sc_hd__or4_4
XFILLER_0_19_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_74_566 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4885_ _4885_/A _4885_/B vssd2 vssd2 vccd2 vccd2 _4887_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_257 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7673_ _7802_/CLK _7673_/D vssd2 vssd2 vccd2 vccd2 _7673_/Q sky130_fd_sc_hd__dfxtp_1
X_6624_ _6551_/A _6551_/B _6546_/X vssd2 vssd2 vccd2 vccd2 _6627_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__5906__B1 _6634_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_15_600 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3836_ _4458_/D _4144_/C vssd2 vssd2 vccd2 vccd2 _4326_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_104_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6555_ _6556_/A _6556_/B vssd2 vssd2 vccd2 vccd2 _6555_/X sky130_fd_sc_hd__and2_1
XFILLER_0_6_387 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5506_ _5506_/A _5506_/B vssd2 vssd2 vccd2 vccd2 _5507_/B sky130_fd_sc_hd__and2_1
X_6486_ _6486_/A _6486_/B vssd2 vssd2 vccd2 vccd2 _6488_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_42_496 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_100_513 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5437_ _5437_/A _5437_/B vssd2 vssd2 vccd2 vccd2 _5439_/B sky130_fd_sc_hd__xnor2_1
X_5368_ _5475_/A _5368_/B vssd2 vssd2 vccd2 vccd2 _5370_/C sky130_fd_sc_hd__and2_1
X_7107_ _7107_/A _7107_/B vssd2 vssd2 vccd2 vccd2 _7109_/B sky130_fd_sc_hd__xor2_1
X_5299_ _5300_/B _5300_/A vssd2 vssd2 vccd2 vccd2 _5299_/X sky130_fd_sc_hd__and2b_1
X_4319_ _4598_/A _4319_/B _4782_/B vssd2 vssd2 vccd2 vccd2 _4367_/B sky130_fd_sc_hd__or3_1
XANTENNA__7080__A _7082_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7038_ _7037_/A _7253_/C _7037_/C vssd2 vssd2 vccd2 vccd2 _7039_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_305 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4209__A _4807_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_349 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_500 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1025 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6424__A _6424_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_77_393 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1069 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_80_514 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_107_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6570__B1 _7045_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5373__B2 _5222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5373__A1 _5374_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7255__A _7291_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_33_452 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4598__B _5374_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_20_146 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_809 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5222__B _5374_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4119__A _4882_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4939__A1 _5210_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4939__B2 _5210_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_68_360 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_56_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_56_511 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_28_224 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1592 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_555 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_83_385 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_71_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4670_ _4670_/A _4670_/B vssd2 vssd2 vccd2 vccd2 _4672_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__5892__B _6812_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_71_558 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_43_249 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_113_137 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6340_ _6783_/A _7037_/A vssd2 vssd2 vccd2 vccd2 _6345_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_3_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_51_271 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_11_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_24_496 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6271_ _6271_/A _6271_/B vssd2 vssd2 vccd2 vccd2 _6272_/B sky130_fd_sc_hd__xnor2_2
X_5222_ _5222_/A _5374_/B vssd2 vssd2 vccd2 vccd2 _5224_/B sky130_fd_sc_hd__nor2_1
X_5153_ _5153_/A vssd2 vssd2 vccd2 vccd2 _5153_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_62 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4104_ _4268_/A _3993_/D _4081_/C _4102_/X _4103_/Y vssd2 vssd2 vccd2 vccd2 _4104_/X
+ sky130_fd_sc_hd__a32o_1
X_5084_ _5084_/A _5084_/B vssd2 vssd2 vccd2 vccd2 _5087_/A sky130_fd_sc_hd__xnor2_1
X_4035_ _7764_/Q _4033_/C _4030_/X _4032_/X _4034_/X vssd2 vssd2 vccd2 vccd2 _4035_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_93_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5986_ _6092_/A _6783_/A vssd2 vssd2 vccd2 vccd2 _5998_/A sky130_fd_sc_hd__nor2_1
XPHY_119 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_108 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_93_149 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4937_ _5042_/A _5550_/A vssd2 vssd2 vccd2 vccd2 _4938_/B sky130_fd_sc_hd__or2_1
XFILLER_0_59_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7725_ _7750_/CLK _7725_/D vssd2 vssd2 vccd2 vccd2 _7725_/Q sky130_fd_sc_hd__dfxtp_1
X_4868_ _5042_/B _5276_/A vssd2 vssd2 vccd2 vccd2 _4869_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_74_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7656_ _7768_/CLK _7656_/D vssd2 vssd2 vccd2 vccd2 _7656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6607_ _6607_/A _6607_/B vssd2 vssd2 vccd2 vccd2 _6608_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_105_627 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3819_ _7803_/Q _3819_/B vssd2 vssd2 vccd2 vccd2 _4522_/C sky130_fd_sc_hd__xor2_4
XANTENNA__6552__B1 _7143_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7587_ _7590_/A vssd2 vssd2 vccd2 vccd2 _7587_/Y sky130_fd_sc_hd__inv_2
X_4799_ _4799_/A _4799_/B vssd2 vssd2 vccd2 vccd2 _4801_/A sky130_fd_sc_hd__xnor2_1
X_6538_ _6538_/A _6615_/B vssd2 vssd2 vccd2 vccd2 _6618_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_30_400 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6469_ _6335_/A _6334_/B _6412_/B _6411_/B _6411_/A vssd2 vssd2 vccd2 vccd2 _6533_/A
+ sky130_fd_sc_hd__a32oi_4
XFILLER_0_42_293 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_100_321 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xoutput160 _7699_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[4] sky130_fd_sc_hd__buf_12
XFILLER_0_100_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6138__B _6973_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6083__A2 _6571_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5042__B _5042_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_108_421 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_53_525 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_53_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_80_333 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4849__A_N _4769_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_80_377 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__5897__A2 _6588_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_21_444 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_33_293 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_103_181 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_606 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_17_32 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_17_65 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5282__B1 _5498_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_88_488 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5840_ _6194_/B _5830_/X _5836_/X _5839_/X vssd2 vssd2 vccd2 vccd2 _5840_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_48_319 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_29_500 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_75_149 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5771_ _6283_/A _5755_/C _5739_/Y _6510_/A vssd2 vssd2 vccd2 vccd2 _5772_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_33_64 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4722_ _4722_/A _4722_/B vssd2 vssd2 vccd2 vccd2 _4757_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_300 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7510_ _7565_/A vssd2 vssd2 vccd2 vccd2 _7510_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_83_193 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_56_385 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7441_ hold127/X _7689_/Q _7451_/S vssd2 vssd2 vccd2 vccd2 _7441_/X sky130_fd_sc_hd__mux2_1
Xinput40 input40/A vssd2 vssd2 vccd2 vccd2 input40/X sky130_fd_sc_hd__clkbuf_1
X_4653_ _4654_/A _4654_/B vssd2 vssd2 vccd2 vccd2 _4653_/Y sky130_fd_sc_hd__nand2_1
X_4584_ _4584_/A _4584_/B vssd2 vssd2 vccd2 vccd2 _4606_/A sky130_fd_sc_hd__xor2_2
Xinput62 wbs_adr_i[20] vssd2 vssd2 vccd2 vccd2 _7340_/B sky130_fd_sc_hd__clkbuf_1
Xinput73 wbs_adr_i[30] vssd2 vssd2 vccd2 vccd2 _7338_/B sky130_fd_sc_hd__clkbuf_1
Xinput51 wbs_adr_i[10] vssd2 vssd2 vccd2 vccd2 _7341_/D sky130_fd_sc_hd__clkbuf_1
X_7372_ _7440_/A _7372_/B vssd2 vssd2 vccd2 vccd2 _7656_/D sky130_fd_sc_hd__and2_1
XANTENNA__7045__D _7253_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xinput95 input95/A vssd2 vssd2 vccd2 vccd2 input95/X sky130_fd_sc_hd__clkbuf_1
Xinput84 input84/A vssd2 vssd2 vccd2 vccd2 input84/X sky130_fd_sc_hd__clkbuf_1
X_6323_ _6398_/A _5659_/B _6396_/B _6322_/X vssd2 vssd2 vccd2 vccd2 _6323_/X sky130_fd_sc_hd__a31o_1
XANTENNA__7623__A _7627_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6254_ _6398_/A _6016_/B _6071_/B _6017_/B _6397_/A vssd2 vssd2 vccd2 vccd2 _6254_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4966__B _5374_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5205_ _5328_/A _5404_/A _5414_/A _5498_/A vssd2 vssd2 vccd2 vccd2 _5206_/B sky130_fd_sc_hd__or4_1
X_6185_ _6185_/A _6185_/B vssd2 vssd2 vccd2 vccd2 _6186_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_94 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_42_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5136_ _5093_/A _5093_/B _5090_/X vssd2 vssd2 vccd2 vccd2 _5139_/A sky130_fd_sc_hd__a21o_1
X_5067_ _5067_/A _5067_/B vssd2 vssd2 vccd2 vccd2 _5128_/B sky130_fd_sc_hd__xor2_4
XANTENNA__4076__A1 _7766_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4018_ _4018_/A _4018_/B _4036_/B vssd2 vssd2 vccd2 vccd2 _4018_/X sky130_fd_sc_hd__and3_1
XFILLER_0_66_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5969_ _5969_/A _5969_/B vssd2 vssd2 vccd2 vccd2 _6068_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_190 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7708_ _7787_/CLK _7708_/D vssd2 vssd2 vccd2 vccd2 _7708_/Q sky130_fd_sc_hd__dfxtp_1
X_7639_ _7641_/A vssd2 vssd2 vccd2 vccd2 _7639_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_62_399 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_62_377 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_50_539 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_50_528 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_105_479 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_30_285 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_100_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4892__A _4962_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_54_19 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_85_458 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_85_447 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5567__A1 _5458_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4116__B _5042_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_108_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_65_193 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_65_182 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_65_160 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_80_130 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_79_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_111_405 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold109 _7444_/X vssd2 vssd2 vccd2 vccd2 _7690_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_104_490 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_95_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_414 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_285 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_425 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5898__A _6283_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4058__A1 _4162_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4058__B2 _7768_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6506__B _7045_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6941_ _6221_/X _6223_/X _7143_/B _6152_/B vssd2 vssd2 vccd2 vccd2 _6944_/A sky130_fd_sc_hd__o211a_1
X_6872_ _6424_/A _6424_/B _6669_/X _7313_/B _6664_/A vssd2 vssd2 vccd2 vccd2 _6872_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_44_74 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_76_469 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5823_ _7807_/D _7336_/A _5865_/A _5818_/Y vssd2 vssd2 vccd2 vccd2 _5824_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_91_417 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_44_322 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_44_300 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5754_ _5748_/X _5749_/Y _5750_/X _5753_/X vssd2 vssd2 vccd2 vccd2 _5760_/B sky130_fd_sc_hd__a211o_1
X_4705_ _4703_/X _4705_/B vssd2 vssd2 vccd2 vccd2 _4709_/A sky130_fd_sc_hd__and2b_1
XANTENNA__4781__A2 _5099_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_72_675 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_72_653 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5685_ _5694_/A _5694_/B _5694_/C _5684_/X _5735_/B vssd2 vssd2 vccd2 vccd2 _5690_/B
+ sky130_fd_sc_hd__o41a_4
XANTENNA__6879__D _7291_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_114_221 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4636_ _4636_/A _4636_/B vssd2 vssd2 vccd2 vccd2 _4639_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_185 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_71_163 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7424_ _7436_/A _7424_/B vssd2 vssd2 vccd2 vccd2 _7680_/D sky130_fd_sc_hd__and2_1
XANTENNA_fanout213_A _6404_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_114_265 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold610 _7814_/Q vssd2 vssd2 vccd2 vccd2 hold610/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 hold621/A vssd2 vssd2 vccd2 vccd2 hold621/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_485 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7355_ hold175/X _7760_/D _7383_/S vssd2 vssd2 vccd2 vccd2 _7355_/X sky130_fd_sc_hd__mux2_1
Xhold643 hold643/A vssd2 vssd2 vccd2 vccd2 hold643/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold632 _7837_/Q vssd2 vssd2 vccd2 vccd2 hold632/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 _7829_/Q vssd2 vssd2 vccd2 vccd2 hold654/X sky130_fd_sc_hd__dlygate4sd3_1
X_6306_ _6306_/A _6306_/B vssd2 vssd2 vccd2 vccd2 _6307_/B sky130_fd_sc_hd__xor2_2
X_4567_ _4898_/A _5276_/A _4498_/B _4497_/B vssd2 vssd2 vccd2 vccd2 _4569_/B sky130_fd_sc_hd__o31a_1
XANTENNA__3881__A _7765_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold665 hold665/A vssd2 vssd2 vccd2 vccd2 hold665/X sky130_fd_sc_hd__dlygate4sd3_1
X_7286_ _7310_/C _7286_/B vssd2 vssd2 vccd2 vccd2 _7833_/D sky130_fd_sc_hd__xnor2_1
X_4498_ _4498_/A _4498_/B vssd2 vssd2 vccd2 vccd2 _4500_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_296 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold687 _7676_/Q vssd2 vssd2 vccd2 vccd2 hold687/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 _3982_/B vssd2 vssd2 vccd2 vccd2 hold676/X sky130_fd_sc_hd__dlygate4sd3_1
X_6237_ _6237_/A _6237_/B vssd2 vssd2 vccd2 vccd2 _6238_/B sky130_fd_sc_hd__xor2_2
Xhold698 _7803_/Q vssd2 vssd2 vccd2 vccd2 _3821_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6168_ _6168_/A _6168_/B vssd2 vssd2 vccd2 vccd2 _6169_/B sky130_fd_sc_hd__xnor2_2
XTAP_970 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_528 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_85_81 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5119_ _5119_/A _5119_/B vssd2 vssd2 vccd2 vccd2 _5122_/A sky130_fd_sc_hd__xnor2_4
XTAP_992 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6099_ _6157_/A _6283_/B vssd2 vssd2 vccd2 vccd2 _6099_/X sky130_fd_sc_hd__and2_1
XANTENNA__6416__B _6973_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5797__B2 _7842_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_67_414 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_94_233 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_67_447 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_39_138 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_94_277 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_35_377 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7226__B2 _7143_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7226__A1 _7145_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6326__B _7181_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5788__A1 _5778_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_98_572 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_81_39 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_58_425 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_105_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_58_458 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_14_44 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6201__A2 _6571_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_73_417 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7438__A _7440_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6342__A _6939_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_26_300 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4212__A1 _7768_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_53_130 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_26_344 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5470_ _5470_/A _5470_/B vssd2 vssd2 vccd2 vccd2 _5472_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_100_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4421_ _4420_/A _4420_/B _4422_/A vssd2 vssd2 vccd2 vccd2 _4480_/B sky130_fd_sc_hd__a21o_1
XANTENNA__6996__B _7181_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_22_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_111_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7140_ _7140_/A _7255_/B vssd2 vssd2 vccd2 vccd2 _7141_/B sky130_fd_sc_hd__nor2_1
X_4352_ _4352_/A _4352_/B vssd2 vssd2 vccd2 vccd2 _4355_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_22_594 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_39_30 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7071_ _6989_/A _7291_/B _7123_/A _7070_/X vssd2 vssd2 vccd2 vccd2 _7072_/B sky130_fd_sc_hd__o22a_1
X_4283_ _4283_/A _4283_/B vssd2 vssd2 vccd2 vccd2 _4285_/B sky130_fd_sc_hd__xnor2_2
XTAP_233 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6022_ _6020_/X _6021_/X _5811_/B vssd2 vssd2 vccd2 vccd2 _6571_/A sky130_fd_sc_hd__o21a_4
XTAP_299 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5779__B2 _7842_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6924_ _6925_/A _6925_/B vssd2 vssd2 vccd2 vccd2 _6924_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_76_244 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6855_ _6855_/A _7255_/B vssd2 vssd2 vccd2 vccd2 _6856_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_9_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_91_225 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6786_ _7047_/A _7094_/A _7143_/A _7143_/B vssd2 vssd2 vccd2 vccd2 _6788_/B sky130_fd_sc_hd__and4_1
X_5806_ _5798_/Y _5800_/Y _5805_/Y _5648_/B vssd2 vssd2 vccd2 vccd2 _5816_/A sky130_fd_sc_hd__a31o_4
X_3998_ _4656_/B _4522_/C _5458_/A vssd2 vssd2 vccd2 vccd2 _4328_/B sky130_fd_sc_hd__and3_1
X_5737_ _6152_/B _5944_/B vssd2 vssd2 vccd2 vccd2 _5737_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_44_174 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7407_ _7452_/A _7407_/B vssd2 vssd2 vccd2 vccd2 _7672_/D sky130_fd_sc_hd__and2_1
X_5668_ _5600_/X _5623_/X _5624_/X _7855_/Q vssd2 vssd2 vccd2 vccd2 _5674_/C sky130_fd_sc_hd__o31a_1
X_4619_ _4619_/A _4619_/B _4619_/C vssd2 vssd2 vccd2 vccd2 _4621_/A sky130_fd_sc_hd__nand3_2
X_5599_ _7842_/Q _5599_/B _5659_/B vssd2 vssd2 vccd2 vccd2 _5599_/X sky130_fd_sc_hd__and3_1
Xhold440 la_data_in[39] vssd2 vssd2 vccd2 vccd2 hold9/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 hold20/X vssd2 vssd2 vccd2 vccd2 _7843_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 input48/X vssd2 vssd2 vccd2 vccd2 hold36/A sky130_fd_sc_hd__dlygate4sd3_1
X_7338_ _7338_/A _7338_/B input70/X input71/X vssd2 vssd2 vccd2 vccd2 _7346_/A sky130_fd_sc_hd__or4bb_1
X_7269_ _7270_/A _7270_/B vssd2 vssd2 vccd2 vccd2 _7303_/A sky130_fd_sc_hd__nor2_1
Xhold495 hold62/X vssd2 vssd2 vccd2 vccd2 _7849_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 la_data_in[14] vssd2 vssd2 vccd2 vccd2 hold21/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 hold41/X vssd2 vssd2 vccd2 vccd2 input10/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5315__B _5315_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5467__B1 _5550_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6427__A _6738_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6431__A2 _5816_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_67_288 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_130 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_63_483 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_152 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7838_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7143__D _7313_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_92_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_25_32 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4433__A1 _5042_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4433__B2 _4863_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4970_ _4970_/A _4970_/B vssd2 vssd2 vccd2 vccd2 _4973_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_86_553 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3921_ _3954_/C _3910_/B _3910_/C _4050_/B vssd2 vssd2 vccd2 vccd2 _3922_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_86_597 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_73_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6640_ _6641_/A _6641_/B vssd2 vssd2 vccd2 vccd2 _6640_/Y sky130_fd_sc_hd__nand2_1
X_3852_ _7793_/Q _7792_/Q _7791_/Q _3888_/B vssd2 vssd2 vccd2 vccd2 _3854_/B sky130_fd_sc_hd__o31a_2
XFILLER_0_41_31 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6571_ _6571_/A _6571_/B _6571_/C _7094_/A vssd2 vssd2 vccd2 vccd2 _6572_/D sky130_fd_sc_hd__and4_1
XFILLER_0_54_450 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5522_ _5561_/A _5561_/B _5522_/C vssd2 vssd2 vccd2 vccd2 _5523_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_26_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_41_86 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7135__B1 _7034_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_41_122 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_112_533 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5453_ _5453_/A _5453_/B vssd2 vssd2 vccd2 vccd2 _5456_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_166 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7334__C _7334_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4404_ _4404_/A _4404_/B vssd2 vssd2 vccd2 vccd2 _4405_/B sky130_fd_sc_hd__xor2_4
X_5384_ _5385_/A _5385_/B vssd2 vssd2 vccd2 vccd2 _5384_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_520 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7123_ _7123_/A _7123_/B vssd2 vssd2 vccd2 vccd2 _7125_/C sky130_fd_sc_hd__xor2_1
X_4335_ _4863_/A _4662_/B _4336_/C vssd2 vssd2 vccd2 vccd2 _4337_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_5_20 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_10_564 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7631__A _7641_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout227 _4880_/B vssd2 vssd2 vccd2 vccd2 _5468_/A sky130_fd_sc_hd__buf_4
Xfanout216 _5105_/B vssd2 vssd2 vccd2 vccd2 _5528_/A sky130_fd_sc_hd__buf_4
X_7054_ _7054_/A _7054_/B vssd2 vssd2 vccd2 vccd2 _7057_/A sky130_fd_sc_hd__xnor2_1
Xfanout249 _3824_/X vssd2 vssd2 vccd2 vccd2 _4809_/B sky130_fd_sc_hd__clkbuf_4
X_4266_ _4264_/Y _4265_/X _5458_/A vssd2 vssd2 vccd2 vccd2 _4266_/X sky130_fd_sc_hd__o21a_1
X_6005_ _5955_/Y _5960_/A _6003_/Y _6004_/X vssd2 vssd2 vccd2 vccd2 _6005_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_66_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4197_ _5548_/A _4305_/A vssd2 vssd2 vccd2 vccd2 _4248_/A sky130_fd_sc_hd__nor2_1
XANTENNA_fanout280_A _7450_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6413__A2 _7037_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_89_391 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1229 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_233 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6907_ _6768_/A _6768_/B _6841_/A _6906_/Y vssd2 vssd2 vccd2 vccd2 _6908_/B sky130_fd_sc_hd__a31o_1
X_6838_ _6838_/A _6838_/B vssd2 vssd2 vccd2 vccd2 _6841_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_49_288 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_9_330 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_107_305 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_18_642 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_107_349 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6769_ _6769_/A _6769_/B _6769_/C vssd2 vssd2 vccd2 vccd2 _7033_/A sky130_fd_sc_hd__and3_1
XFILLER_0_60_442 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6710__A _7047_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_60_497 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_32_188 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
Xhold270 hold270/A vssd2 vssd2 vccd2 vccd2 la_data_out[2] sky130_fd_sc_hd__buf_12
Xhold281 hold634/X vssd2 vssd2 vccd2 vccd2 hold635/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 hold292/A vssd2 vssd2 vccd2 vccd2 la_data_out[14] sky130_fd_sc_hd__buf_12
XANTENNA__4884__B _5030_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_99_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6157__A _6157_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_317 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_68_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_28_406 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_55_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7138__D _7253_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_70_228 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_23_100 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_36_483 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_11_306 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__3963__B _4050_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_23_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_87_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_23_199 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4140__A _4807_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4120_ _4656_/A _5030_/A vssd2 vssd2 vccd2 vccd2 _4120_/X sky130_fd_sc_hd__and2_1
X_4051_ _7727_/D _5455_/A vssd2 vssd2 vccd2 vccd2 _4052_/B sky130_fd_sc_hd__nand2_1
Xinput5 input5/A vssd2 vssd2 vccd2 vccd2 input5/X sky130_fd_sc_hd__buf_1
XFILLER_0_36_64 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7810_ _7814_/CLK _7810_/D _7569_/Y vssd2 vssd2 vccd2 vccd2 _7810_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_520 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_59_575 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4953_ _5029_/A _5105_/B _5550_/B _4882_/A vssd2 vssd2 vccd2 vccd2 _4956_/A sky130_fd_sc_hd__o22ai_1
X_7741_ _7787_/CLK _7741_/D _7500_/Y vssd2 vssd2 vccd2 vccd2 _7741_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_394 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7672_ _7768_/CLK _7672_/D vssd2 vssd2 vccd2 vccd2 _7672_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6159__A1 _6282_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4315__A _4809_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3904_ _3904_/A _3904_/B _3904_/C vssd2 vssd2 vccd2 vccd2 _4708_/A sky130_fd_sc_hd__and3_4
X_6623_ _6564_/A _6564_/B _6567_/A vssd2 vssd2 vccd2 vccd2 _6627_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_52_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4884_ _5030_/A _5030_/B _5326_/A vssd2 vssd2 vccd2 vccd2 _4885_/B sky130_fd_sc_hd__and3_1
XFILLER_0_74_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3835_ _7800_/Q _3835_/B vssd2 vssd2 vccd2 vccd2 _4006_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_461 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__7626__A _7627_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6554_ _6556_/A _6556_/B vssd2 vssd2 vccd2 vccd2 _6554_/X sky130_fd_sc_hd__or2_1
X_6485_ _6486_/A _6486_/B vssd2 vssd2 vccd2 vccd2 _6566_/A sky130_fd_sc_hd__and2b_1
XANTENNA__4590__B1 _5222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5505_ _5506_/A _5506_/B vssd2 vssd2 vccd2 vccd2 _5539_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_72_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5436_ _5480_/B _5436_/B _5437_/B vssd2 vssd2 vccd2 vccd2 _5486_/A sky130_fd_sc_hd__or3_1
XFILLER_0_112_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_10_372 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5367_ _5366_/A _5498_/D _5366_/C vssd2 vssd2 vccd2 vccd2 _5368_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_93 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5298_ _5240_/A _5240_/B _5238_/X vssd2 vssd2 vccd2 vccd2 _5300_/B sky130_fd_sc_hd__a21oi_2
X_7106_ _7106_/A _7106_/B vssd2 vssd2 vccd2 vccd2 _7107_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_10_394 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4318_ _4314_/X _4317_/X _4214_/B vssd2 vssd2 vccd2 vccd2 _4318_/Y sky130_fd_sc_hd__o21ai_2
X_7037_ _7037_/A _7253_/C _7037_/C vssd2 vssd2 vccd2 vccd2 _7153_/A sky130_fd_sc_hd__or3_2
X_4249_ _4893_/A _4020_/B _4122_/D _7766_/Q _4815_/B vssd2 vssd2 vccd2 vccd2 _4249_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4645__A1 _4810_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_93_81 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_69_317 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4209__B _5042_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6705__A _6783_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1004 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_350 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1037 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_236 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_107_113 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_18_472 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6570__B2 _6973_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_52_228 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__7536__A _7557_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5373__A2 _5468_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7255__B _7255_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6858__C1 _7143_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_57_19 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4895__A _5099_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4119__B _4863_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__4939__A2 _5222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1560 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_567 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_56_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_28_236 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_113_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_56_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_43_206 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_98_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6350__A _6664_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7446__A _7452_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_113_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_24_464 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_113_149 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6270_ _6271_/B _6271_/A vssd2 vssd2 vccd2 vccd2 _6270_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_51_294 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7181__A _7181_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5221_ _4266_/X _4270_/X _4814_/Y _3996_/B vssd2 vssd2 vccd2 vccd2 _5224_/A sky130_fd_sc_hd__o211a_1
X_5152_ _5276_/A _5315_/B _5154_/A vssd2 vssd2 vccd2 vccd2 _5153_/A sky130_fd_sc_hd__or3_1
X_4103_ _4103_/A _4103_/B vssd2 vssd2 vccd2 vccd2 _4103_/Y sky130_fd_sc_hd__nor2_1
X_5083_ _5366_/A _5431_/A vssd2 vssd2 vccd2 vccd2 _5084_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_47_74 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4627__A1 _4268_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_2_10 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4034_ _4315_/B _4070_/D _4034_/C vssd2 vssd2 vccd2 vccd2 _4034_/X sky130_fd_sc_hd__and3_1
XFILLER_0_66_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5985_ _5985_/A _5985_/B vssd2 vssd2 vccd2 vccd2 _6003_/A sky130_fd_sc_hd__xor2_1
XPHY_109 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_47_512 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7724_ _7750_/CLK _7724_/D vssd2 vssd2 vccd2 vccd2 _7724_/Q sky130_fd_sc_hd__dfxtp_1
X_4936_ _4938_/A vssd2 vssd2 vccd2 vccd2 _4936_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7329__B1 _6669_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_19_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_19_236 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_19_247 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4867_ _4865_/X _4867_/B vssd2 vssd2 vccd2 vccd2 _4869_/A sky130_fd_sc_hd__and2b_1
X_7655_ _7802_/CLK _7655_/D vssd2 vssd2 vccd2 vccd2 _7655_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_10 wbs_adr_i[2] vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_19_258 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6606_ _6607_/A _6607_/B vssd2 vssd2 vccd2 vccd2 _6606_/Y sky130_fd_sc_hd__nor2_1
X_7586_ _7590_/A vssd2 vssd2 vccd2 vccd2 _7586_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_62_537 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7356__A _7436_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3818_ _7804_/Q _3818_/B vssd2 vssd2 vccd2 vccd2 _4656_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_34_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6537_ _6537_/A _6537_/B vssd2 vssd2 vccd2 vccd2 _6615_/B sky130_fd_sc_hd__xor2_2
XANTENNA__4563__B1 _4782_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4798_ _4882_/A _5105_/B _4799_/A vssd2 vssd2 vccd2 vccd2 _4798_/X sky130_fd_sc_hd__or3_1
X_6468_ _6458_/Y _6462_/B _6456_/Y vssd2 vssd2 vccd2 vccd2 _6538_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_100_333 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6399_ _6396_/Y _6397_/Y _6398_/Y _5653_/C vssd2 vssd2 vccd2 vccd2 _7222_/A sky130_fd_sc_hd__a31oi_4
Xoutput161 _7700_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[5] sky130_fd_sc_hd__buf_12
Xoutput150 _7719_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[24] sky130_fd_sc_hd__buf_12
X_5419_ _5420_/B _5421_/B vssd2 vssd2 vccd2 vccd2 _5472_/A sky130_fd_sc_hd__nor2_1
XANTENNA__5042__C _5374_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_103 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_97_467 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_97_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_69_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_69_147 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_38_512 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_84_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6791__A1 _6939_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_108_411 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_53_515 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_108_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_53_537 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__3794__A _4268_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_80_345 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_18_291 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_581 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_250 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_21_456 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_193 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_607 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4857__A1 _4598_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_618 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_401 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_17_44 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5282__B2 _5431_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5282__A1 _5404_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_48_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_8_428 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5770_ _5845_/B _5845_/C vssd2 vssd2 vccd2 vccd2 _5853_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_29_556 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1390 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_109 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4721_ _4722_/A _4722_/B vssd2 vssd2 vccd2 vccd2 _4772_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_29_578 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4652_ _4654_/A _4654_/B vssd2 vssd2 vccd2 vccd2 _4652_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__7176__A _7224_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7440_ _7440_/A _7440_/B vssd2 vssd2 vccd2 vccd2 _7688_/D sky130_fd_sc_hd__and2_1
Xinput30 input30/A vssd2 vssd2 vccd2 vccd2 input30/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__7326__D _7326_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_71_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4583_ _4583_/A _4583_/B vssd2 vssd2 vccd2 vccd2 _4584_/B sky130_fd_sc_hd__xor2_2
Xinput41 input41/A vssd2 vssd2 vccd2 vccd2 input41/X sky130_fd_sc_hd__clkbuf_1
Xinput52 wbs_adr_i[11] vssd2 vssd2 vccd2 vccd2 _7341_/C sky130_fd_sc_hd__clkbuf_1
Xinput63 wbs_adr_i[21] vssd2 vssd2 vccd2 vccd2 _7340_/A sky130_fd_sc_hd__clkbuf_1
X_7371_ hold221/X _7768_/D _7383_/S vssd2 vssd2 vccd2 vccd2 _7372_/B sky130_fd_sc_hd__mux2_1
Xinput85 input85/A vssd2 vssd2 vccd2 vccd2 input85/X sky130_fd_sc_hd__clkbuf_1
Xinput96 input96/A vssd2 vssd2 vccd2 vccd2 input96/X sky130_fd_sc_hd__clkbuf_1
Xinput74 wbs_adr_i[31] vssd2 vssd2 vccd2 vccd2 _7338_/A sky130_fd_sc_hd__clkbuf_1
X_6322_ _6397_/A _5659_/A _6194_/B _6074_/A _7313_/A vssd2 vssd2 vccd2 vccd2 _6322_/X
+ sky130_fd_sc_hd__a32o_1
X_6253_ _6253_/A _6253_/B _6253_/C vssd2 vssd2 vccd2 vccd2 _6253_/X sky130_fd_sc_hd__and3_1
XFILLER_0_110_675 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_58_73 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5204_ _5404_/A _5414_/A _5498_/A _5328_/A vssd2 vssd2 vccd2 vccd2 _5206_/A sky130_fd_sc_hd__o22ai_1
X_6184_ _6184_/A _6184_/B _6185_/A vssd2 vssd2 vccd2 vccd2 _6184_/X sky130_fd_sc_hd__or3_1
X_5135_ _5123_/A _5123_/B _5121_/X vssd2 vssd2 vccd2 vccd2 _5195_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_35_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_98_209 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5066_ _5067_/A _5067_/B vssd2 vssd2 vccd2 vccd2 _5250_/A sky130_fd_sc_hd__and2_1
X_4017_ _4017_/A _4017_/B vssd2 vssd2 vccd2 vccd2 _4779_/A sky130_fd_sc_hd__and2_2
XFILLER_0_94_415 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_94_448 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5968_ _5968_/A _5969_/B vssd2 vssd2 vccd2 vccd2 _5968_/X sky130_fd_sc_hd__or2_1
XANTENNA__6773__A1 _6707_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_47_331 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4919_ _4919_/A _4919_/B vssd2 vssd2 vccd2 vccd2 _4920_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_81_109 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_75_673 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7707_ _7787_/CLK _7707_/D vssd2 vssd2 vccd2 vccd2 _7707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_515 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_47_397 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5899_ _7847_/Q _5937_/B _5935_/D _6158_/A vssd2 vssd2 vccd2 vccd2 _5899_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_35_537 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_548 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_7_461 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7638_ _7641_/A vssd2 vssd2 vccd2 vccd2 _7638_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_105_436 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7569_ _7613_/A vssd2 vssd2 vccd2 vccd2 _7569_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_50_518 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_15_294 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_30_242 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_100_141 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_58_607 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_57_106 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_57_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5567__A2 _5431_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_72_109 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_38_342 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_93_492 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5972__C1 _5736_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_26_515 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_26_548 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_81_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_79_39 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4527__B1 _4965_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_13_209 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_111_417 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_21_264 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_95_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_415 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5898__B _5992_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6940_ _6940_/A _6940_/B vssd2 vssd2 vccd2 vccd2 _6950_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_253 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6871_ _6871_/A _6871_/B vssd2 vssd2 vccd2 vccd2 _6891_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__3927__C_N _4050_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5822_ _5818_/Y _5865_/A _7336_/A _7807_/D vssd2 vssd2 vccd2 vccd2 _5824_/A sky130_fd_sc_hd__o211ai_1
XANTENNA__6803__A _7037_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5753_ _7841_/Q _6283_/B _6358_/B vssd2 vssd2 vccd2 vccd2 _5753_/X sky130_fd_sc_hd__and3_1
XFILLER_0_84_492 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4704_ _4779_/A _4704_/B _5142_/C _5076_/D vssd2 vssd2 vccd2 vccd2 _4705_/B sky130_fd_sc_hd__or4_1
XFILLER_0_60_52 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_60_41 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_56_161 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_29_375 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_44_334 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5684_ _7879_/Q _7880_/Q vssd2 vssd2 vccd2 vccd2 _5684_/X sky130_fd_sc_hd__or2_1
X_4635_ _4633_/X _4635_/B vssd2 vssd2 vccd2 vccd2 _4636_/B sky130_fd_sc_hd__and2b_1
XANTENNA__7180__A1 _7051_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7423_ hold175/X _7680_/Q _7451_/S vssd2 vssd2 vccd2 vccd2 _7423_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_518 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_114_277 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xhold611 hold611/A vssd2 vssd2 vccd2 vccd2 hold611/X sky130_fd_sc_hd__dlygate4sd3_1
X_4566_ _4566_/A _4566_/B vssd2 vssd2 vccd2 vccd2 _4569_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__7180__B2 _6479_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_fanout206_A _5011_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7354_ _7436_/A _7354_/B vssd2 vssd2 vccd2 vccd2 _7647_/D sky130_fd_sc_hd__and2_1
Xhold600 la_data_in[0] vssd2 vssd2 vccd2 vccd2 hold95/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7634__A _7641_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold633 hold633/A vssd2 vssd2 vccd2 vccd2 hold633/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 _7827_/Q vssd2 vssd2 vccd2 vccd2 hold644/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_439 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6305_ _6306_/A _6306_/B vssd2 vssd2 vccd2 vccd2 _6305_/Y sky130_fd_sc_hd__nor2_1
Xhold622 _7809_/Q vssd2 vssd2 vccd2 vccd2 hold622/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_72 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
Xhold655 hold655/A vssd2 vssd2 vccd2 vccd2 hold655/X sky130_fd_sc_hd__dlygate4sd3_1
X_7285_ _7310_/A _7219_/B _7310_/B _7336_/A vssd2 vssd2 vccd2 vccd2 _7286_/B sky130_fd_sc_hd__o31ai_1
Xhold666 _7818_/Q vssd2 vssd2 vccd2 vccd2 hold666/X sky130_fd_sc_hd__dlygate4sd3_1
X_4497_ _4497_/A _4497_/B vssd2 vssd2 vccd2 vccd2 _4498_/B sky130_fd_sc_hd__nand2_1
Xhold688 _7666_/Q vssd2 vssd2 vccd2 vccd2 hold688/X sky130_fd_sc_hd__dlygate4sd3_1
X_6236_ _6237_/A _6237_/B vssd2 vssd2 vccd2 vccd2 _6236_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7483__A2 _7483_/A2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold699 _3821_/X vssd2 vssd2 vccd2 vccd2 _3822_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6167_ _6168_/B _6168_/A vssd2 vssd2 vccd2 vccd2 _6167_/Y sky130_fd_sc_hd__nand2b_1
XTAP_960 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5118_ _5118_/A _5118_/B vssd2 vssd2 vccd2 vccd2 _5119_/B sky130_fd_sc_hd__xor2_4
XTAP_993 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6098_ _6510_/A _5935_/X _6096_/Y _6097_/X vssd2 vssd2 vccd2 vccd2 _6098_/X sky130_fd_sc_hd__a211o_1
XANTENNA__6416__C _6989_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5049_ _4974_/A _4974_/B _4972_/Y vssd2 vssd2 vccd2 vccd2 _5051_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_79_275 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_39_117 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_94_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6713__A _6939_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_94_289 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_63_610 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_35_356 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_63_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__3980__A1 _7761_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_23_518 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_62_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7474__A2 _7483_/A2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7226__A2 _7313_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5788__A2 _5786_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_85_212 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_105_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_14_56 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_651 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6342__B _6973_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_73_429 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_66_470 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_39_673 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_30_22 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4143__A _7768_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_81_473 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_54_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_14_518 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4420_ _4420_/A _4420_/B vssd2 vssd2 vccd2 vccd2 _4422_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_111_225 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4351_ _4351_/A _4351_/B vssd2 vssd2 vccd2 vccd2 _4352_/B sky130_fd_sc_hd__xnor2_2
X_7070_ _7070_/A _7070_/B _7070_/C vssd2 vssd2 vccd2 vccd2 _7070_/X sky130_fd_sc_hd__and3_1
X_4282_ _4044_/A _4044_/B _4966_/A vssd2 vssd2 vccd2 vccd2 _4283_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__7465__A2 _7454_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_39_75 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XTAP_256 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6021_ _6397_/A _5825_/X _6015_/X _6017_/X _6019_/X vssd2 vssd2 vccd2 vccd2 _6021_/X
+ sky130_fd_sc_hd__a2111o_2
XTAP_289 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5779__A2 _6588_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6923_ _7037_/A _7224_/A vssd2 vssd2 vccd2 vccd2 _6925_/B sky130_fd_sc_hd__or2_1
XFILLER_0_49_426 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7629__A _7629_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6854_ _6854_/A _6854_/B vssd2 vssd2 vccd2 vccd2 _6856_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_237 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_57_481 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6785_ _7094_/A _7143_/A _7143_/B _7047_/A vssd2 vssd2 vccd2 vccd2 _6785_/X sky130_fd_sc_hd__a22o_1
XANTENNA__7348__B _7436_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3997_ _4457_/B _4458_/C vssd2 vssd2 vccd2 vccd2 _4380_/B sky130_fd_sc_hd__nor2_1
X_5805_ _5803_/X _5804_/X _6253_/C vssd2 vssd2 vccd2 vccd2 _5805_/Y sky130_fd_sc_hd__o21ai_1
X_5736_ _7872_/Q _5736_/B vssd2 vssd2 vccd2 vccd2 _5736_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_60_613 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_45_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_17_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5667_ _7855_/Q _5661_/B _5658_/Y _5666_/X _5664_/X vssd2 vssd2 vccd2 vccd2 _5667_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_44_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7406_ hold221/X _7784_/D _7418_/S vssd2 vssd2 vccd2 vccd2 _7407_/B sky130_fd_sc_hd__mux2_1
XANTENNA__7364__A _7440_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_32_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_32_348 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4618_ _4618_/A _4618_/B vssd2 vssd2 vccd2 vccd2 _4619_/C sky130_fd_sc_hd__xnor2_2
X_5598_ _7867_/Q _5598_/B vssd2 vssd2 vccd2 vccd2 _5653_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_13_540 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_32_359 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold452 la_data_in[46] vssd2 vssd2 vccd2 vccd2 hold25/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 hold9/X vssd2 vssd2 vccd2 vccd2 input33/A sky130_fd_sc_hd__dlygate4sd3_1
X_7337_ _6629_/B _6629_/C _6669_/X _7336_/B _7336_/A vssd2 vssd2 vccd2 vccd2 _7337_/X
+ sky130_fd_sc_hd__a32o_1
Xhold430 input2/X vssd2 vssd2 vccd2 vccd2 hold6/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 hold36/X vssd2 vssd2 vccd2 vccd2 _7880_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4549_ _4479_/A _4480_/A _4479_/B vssd2 vssd2 vccd2 vccd2 _4551_/C sky130_fd_sc_hd__a21o_1
X_7268_ _7300_/A _7268_/B vssd2 vssd2 vccd2 vccd2 _7270_/B sky130_fd_sc_hd__or2_1
Xhold485 hold21/X vssd2 vssd2 vccd2 vccd2 input6/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7456__A2 _7454_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold496 la_data_in[17] vssd2 vssd2 vccd2 vccd2 hold51/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 input10/X vssd2 vssd2 vccd2 vccd2 hold42/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5315__C _5498_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6219_ _5816_/A _5816_/B _7045_/A vssd2 vssd2 vccd2 vccd2 _6228_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__5467__A1 _5498_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5467__B2 _5404_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7199_ _7199_/A _7199_/B _7199_/C vssd2 vssd2 vccd2 vccd2 _7200_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_99_337 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_790 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_55_407 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_95_598 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_82_226 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6162__B _7094_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_48_492 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4898__A _4898_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3953__A1 _4050_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_23_315 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_63_495 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_23_348 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_31_370 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_86_510 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4433__A2 _4711_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3920_ _7763_/Q _4252_/B vssd2 vssd2 vccd2 vccd2 _3920_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_25_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_86_587 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3851_ _7793_/Q _3851_/B vssd2 vssd2 vccd2 vccd2 _4084_/B sky130_fd_sc_hd__xnor2_1
X_6570_ _6571_/B _6571_/C _7045_/A _6973_/A vssd2 vssd2 vccd2 vccd2 _6572_/C sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_73_237 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_41_43 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_109_391 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5521_ _5561_/B _5522_/C _5561_/A vssd2 vssd2 vccd2 vccd2 _5544_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_112_501 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_81_292 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_41_101 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5452_ _5451_/A _5451_/B _5453_/A vssd2 vssd2 vccd2 vccd2 _5488_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_41_145 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_41_156 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_112_545 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4403_ _4404_/A _4404_/B vssd2 vssd2 vccd2 vccd2 _4403_/Y sky130_fd_sc_hd__nor2_1
X_5383_ _5334_/B _5379_/B _5336_/B _5336_/A vssd2 vssd2 vccd2 vccd2 _5385_/B sky130_fd_sc_hd__o22a_2
XFILLER_0_1_220 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_112_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7122_ _7123_/A _7123_/B vssd2 vssd2 vccd2 vccd2 _7169_/B sky130_fd_sc_hd__nand2_1
X_4334_ _4962_/A _4966_/A vssd2 vssd2 vccd2 vccd2 _4336_/C sky130_fd_sc_hd__or2_1
XFILLER_0_22_381 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7053_ _7237_/A _7181_/A vssd2 vssd2 vccd2 vccd2 _7054_/B sky130_fd_sc_hd__nor2_1
Xfanout206 _5011_/A vssd2 vssd2 vccd2 vccd2 _4896_/A sky130_fd_sc_hd__clkbuf_8
Xfanout217 _5145_/B vssd2 vssd2 vccd2 vccd2 _5550_/A sky130_fd_sc_hd__clkbuf_8
X_6004_ _6003_/B _6003_/C _6003_/A vssd2 vssd2 vccd2 vccd2 _6004_/X sky130_fd_sc_hd__a21o_1
X_4265_ _4328_/A _4519_/B _3820_/Y _4745_/A _7767_/Q vssd2 vssd2 vccd2 vccd2 _4265_/X
+ sky130_fd_sc_hd__a32o_1
X_4196_ _4196_/A _4196_/B vssd2 vssd2 vccd2 vccd2 _4305_/A sky130_fd_sc_hd__and2_1
XANTENNA__4121__B2 _7765_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_fanout273_A _7771_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_96_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_89_370 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1219 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_201 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6906_ _6762_/A _6836_/Y _6838_/B vssd2 vssd2 vccd2 vccd2 _6906_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_576 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_77_565 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_49_256 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7886_ _7886_/CLK _7886_/D _7645_/Y vssd2 vssd2 vccd2 vccd2 _7886_/Q sky130_fd_sc_hd__dfrtp_4
X_6837_ _6839_/A _6839_/B vssd2 vssd2 vccd2 vccd2 _6838_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_64_226 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_64_215 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_107_317 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_9_386 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6768_ _6768_/A _6768_/B vssd2 vssd2 vccd2 vccd2 _6909_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_164 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_18_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6699_ _6700_/A _6700_/B vssd2 vssd2 vccd2 vccd2 _6834_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6710__B _7143_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7094__A _7094_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5719_ _5735_/B _7875_/Q _5731_/B vssd2 vssd2 vccd2 vccd2 _5720_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_60_454 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_20_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold271 hold632/X vssd2 vssd2 vccd2 vccd2 hold633/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold260 hold260/A vssd2 vssd2 vccd2 vccd2 la_data_out[6] sky130_fd_sc_hd__buf_12
Xhold293 hold644/X vssd2 vssd2 vccd2 vccd2 hold645/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 hold282/A vssd2 vssd2 vccd2 vccd2 la_data_out[13] sky130_fd_sc_hd__buf_12
XFILLER_0_99_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_87_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__3797__A _4328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_68_587 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_28_418 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_55_237 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_11_24 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_36_473 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_63_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_51_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_635 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_11_79 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_87_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_23_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4140__B _4863_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4050_ _4050_/A _4050_/B vssd2 vssd2 vccd2 vccd2 _5548_/A sky130_fd_sc_hd__xnor2_4
Xinput6 input6/A vssd2 vssd2 vccd2 vccd2 input6/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5851__B2 _7843_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5851__A1 _7845_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_340 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4952_ _4885_/A _4885_/B _4882_/X vssd2 vssd2 vccd2 vccd2 _4959_/B sky130_fd_sc_hd__a21bo_1
X_7740_ _7787_/CLK _7740_/D _7499_/Y vssd2 vssd2 vccd2 vccd2 _7740_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_362 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6514__C _7294_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4883_ _4883_/A _4883_/B vssd2 vssd2 vccd2 vccd2 _4885_/A sky130_fd_sc_hd__xnor2_1
X_7671_ _7802_/CLK _7671_/D vssd2 vssd2 vccd2 vccd2 _7671_/Q sky130_fd_sc_hd__dfxtp_1
X_3903_ _4082_/B _4002_/C _3890_/X _3900_/X wire228/X vssd2 vssd2 vccd2 vccd2 _3904_/C
+ sky130_fd_sc_hd__a311oi_4
X_6622_ _6765_/A _6617_/B _6612_/Y vssd2 vssd2 vccd2 vccd2 _6695_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_237 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3834_ _7800_/Q _3835_/B vssd2 vssd2 vccd2 vccd2 _4144_/C sky130_fd_sc_hd__xor2_4
XFILLER_0_15_613 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_104_309 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6553_ _5991_/X _5993_/X _7143_/A _5781_/B vssd2 vssd2 vccd2 vccd2 _6556_/B sky130_fd_sc_hd__o211a_1
XFILLER_0_42_421 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_27_484 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_495 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6484_ _6402_/A _7145_/A _6406_/B _6405_/B vssd2 vssd2 vccd2 vccd2 _6486_/B sky130_fd_sc_hd__a31o_1
XANTENNA__4590__B2 _4962_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5504_ _5406_/A _5431_/B _5469_/A _5469_/B vssd2 vssd2 vccd2 vccd2 _5506_/B sky130_fd_sc_hd__o22a_1
X_5435_ _5390_/A _5390_/B _5384_/X vssd2 vssd2 vccd2 vccd2 _5437_/B sky130_fd_sc_hd__o21a_1
XANTENNA__4050__B _4050_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_65_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_77_61 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5366_ _5366_/A _5498_/D _5366_/C vssd2 vssd2 vccd2 vccd2 _5475_/A sky130_fd_sc_hd__or3_1
X_7105_ _7106_/A _7106_/B vssd2 vssd2 vccd2 vccd2 _7105_/Y sky130_fd_sc_hd__nor2_1
X_5297_ _5297_/A _5297_/B vssd2 vssd2 vccd2 vccd2 _5300_/A sky130_fd_sc_hd__xnor2_2
X_4317_ _4268_/A _4160_/B _4316_/X _4427_/A _4315_/X vssd2 vssd2 vccd2 vccd2 _4317_/X
+ sky130_fd_sc_hd__a221o_1
X_7036_ _6973_/B _7253_/D _6670_/Y _6973_/A vssd2 vssd2 vccd2 vccd2 _7037_/C sky130_fd_sc_hd__o22a_1
X_4248_ _4248_/A _4305_/B vssd2 vssd2 vccd2 vccd2 _7732_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__4645__A2 _5406_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_93_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7044__B1 _7222_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4179_ _4180_/A _4180_/B vssd2 vssd2 vccd2 vccd2 _4179_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6705__B _6705_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1038 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6424__C _7197_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_92_321 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7869_ _7870_/CLK _7869_/D _7628_/Y vssd2 vssd2 vccd2 vccd2 _7869_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_248 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_107_125 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_92_365 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_107_169 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_80_549 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_45_281 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6858__B1 _6152_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_33_487 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_20_137 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7552__A _7557_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4895__B _5220_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5800__A _6158_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_137 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1550 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_181 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_90 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_113_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6350__B _7047_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_22_78 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_24_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_98_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_36_292 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_24_487 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5220_ _5220_/A _5468_/A vssd2 vssd2 vccd2 vccd2 _5225_/A sky130_fd_sc_hd__or2_1
XANTENNA__7181__B _7253_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5151_ _5276_/A _5315_/B _5154_/A vssd2 vssd2 vccd2 vccd2 _5151_/X sky130_fd_sc_hd__o21a_1
X_5082_ _5082_/A _5082_/B vssd2 vssd2 vccd2 vccd2 _5084_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6077__A1 _7847_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6077__B2 _7848_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4102_ _4002_/A _4002_/B _4002_/C _4101_/Y _4099_/X vssd2 vssd2 vccd2 vccd2 _4102_/X
+ sky130_fd_sc_hd__a41o_1
X_4033_ _7768_/Q _4214_/B _4033_/C vssd2 vssd2 vccd2 vccd2 _4034_/C sky130_fd_sc_hd__and3_1
XFILLER_0_78_126 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_78_148 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_63_74 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4326__A _4656_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5984_ _6550_/A _5984_/B vssd2 vssd2 vccd2 vccd2 _5985_/B sky130_fd_sc_hd__nor2_1
X_7723_ _7723_/CLK _7723_/D vssd2 vssd2 vccd2 vccd2 _7723_/Q sky130_fd_sc_hd__dfxtp_1
X_4935_ _4935_/A _4935_/B vssd2 vssd2 vccd2 vccd2 _4938_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__7329__A1 _6588_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7637__A _7641_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_74_376 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_74_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4866_ _5210_/A _5210_/B _4965_/B _5222_/A vssd2 vssd2 vccd2 vccd2 _4867_/B sky130_fd_sc_hd__or4_1
XFILLER_0_62_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7654_ _7798_/CLK _7654_/D vssd2 vssd2 vccd2 vccd2 _7654_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_11 wbs_dat_i[5] vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_34_207 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6605_ _6528_/A _6528_/B _6526_/Y vssd2 vssd2 vccd2 vccd2 _6607_/B sky130_fd_sc_hd__a21boi_1
X_7585_ _7590_/A vssd2 vssd2 vccd2 vccd2 _7585_/Y sky130_fd_sc_hd__inv_2
X_4797_ wire212/X _4881_/A2 _5528_/A vssd2 vssd2 vccd2 vccd2 _4799_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3817_ _7804_/Q _3818_/B vssd2 vssd2 vccd2 vccd2 _4745_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_27_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6536_ _6536_/A _6536_/B vssd2 vssd2 vccd2 vccd2 _6537_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__4563__B2 _4896_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4563__A1 _4966_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_15_432 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_104_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_100_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6467_ _7336_/A _6467_/B vssd2 vssd2 vccd2 vccd2 _6539_/A sky130_fd_sc_hd__nand2_1
XANTENNA__7372__A _7440_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6398_ _6398_/A _6398_/B vssd2 vssd2 vccd2 vccd2 _6398_/Y sky130_fd_sc_hd__nand2_1
Xoutput140 _7710_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[15] sky130_fd_sc_hd__buf_12
Xoutput151 _7720_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[25] sky130_fd_sc_hd__buf_12
X_5418_ _5461_/B _5418_/B vssd2 vssd2 vccd2 vccd2 _5421_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_100_345 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5349_ _5349_/A _5349_/B vssd2 vssd2 vccd2 vccd2 _5350_/B sky130_fd_sc_hd__nand2_1
Xoutput162 _7701_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[6] sky130_fd_sc_hd__buf_12
XANTENNA__7265__B1 _7224_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7019_ _7019_/A _7019_/B vssd2 vssd2 vccd2 vccd2 _7020_/B sky130_fd_sc_hd__and2_1
XANTENNA__5042__D _5528_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5620__A _7846_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6435__B _7222_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_77_192 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6791__A2 _7181_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_65_376 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_65_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_65_343 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_38_568 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xwire212 _4044_/A vssd2 vssd2 vccd2 vccd2 wire212/X sky130_fd_sc_hd__buf_4
XFILLER_0_92_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_80_357 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_18_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_33_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_110_109 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_61_593 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_161 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4857__A2 _5431_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_608 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_88_413 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5282__A2 _5406_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4146__A _7765_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_671 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_33_11 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1391 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_674 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4720_ _4720_/A _4720_/B vssd2 vssd2 vccd2 vccd2 _4722_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_56_365 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4651_ _4651_/A _4651_/B vssd2 vssd2 vccd2 vccd2 _4654_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__7176__B _7253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xinput31 input31/A vssd2 vssd2 vccd2 vccd2 input31/X sky130_fd_sc_hd__clkbuf_1
Xinput20 input20/A vssd2 vssd2 vccd2 vccd2 input20/X sky130_fd_sc_hd__clkbuf_1
Xinput42 input42/A vssd2 vssd2 vccd2 vccd2 input42/X sky130_fd_sc_hd__clkbuf_1
X_4582_ _4583_/A _4583_/B vssd2 vssd2 vccd2 vccd2 _4582_/Y sky130_fd_sc_hd__nor2_1
X_7370_ _7452_/A _7370_/B vssd2 vssd2 vccd2 vccd2 _7655_/D sky130_fd_sc_hd__and2_1
Xinput53 wbs_adr_i[12] vssd2 vssd2 vccd2 vccd2 _7343_/B sky130_fd_sc_hd__buf_1
Xinput64 input64/A vssd2 vssd2 vccd2 vccd2 _7340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_262 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6321_ _6272_/A _6272_/B _6270_/X vssd2 vssd2 vccd2 vccd2 _6337_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_12_446 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
Xinput75 input75/A vssd2 vssd2 vccd2 vccd2 input75/X sky130_fd_sc_hd__clkbuf_1
Xinput86 input86/A vssd2 vssd2 vccd2 vccd2 input86/X sky130_fd_sc_hd__clkbuf_1
Xinput97 input97/A vssd2 vssd2 vccd2 vccd2 input97/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_178 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_110_632 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6252_ _7850_/Q _7313_/A _6398_/B _6283_/A vssd2 vssd2 vccd2 vccd2 _6252_/X sky130_fd_sc_hd__a22o_1
X_6183_ _6184_/A _6184_/B vssd2 vssd2 vccd2 vccd2 _6185_/B sky130_fd_sc_hd__nor2_1
X_5203_ _5151_/X _5153_/Y _5156_/B _5159_/A vssd2 vssd2 vccd2 vccd2 _5219_/A sky130_fd_sc_hd__o31ai_2
XFILLER_0_58_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5134_ _5455_/A _5357_/A vssd2 vssd2 vccd2 vccd2 _5198_/A sky130_fd_sc_hd__nand2_1
X_5065_ _4990_/A _4990_/B _4988_/Y vssd2 vssd2 vccd2 vccd2 _5067_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_74_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA_fanout186_A _6425_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6470__A1 _5819_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4016_ _4001_/Y _4005_/Y _4014_/X _4015_/Y _3893_/D vssd2 vssd2 vccd2 vccd2 _4017_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_28_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_79_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_66_118 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6222__B2 _6283_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5967_ _5967_/A _5967_/B vssd2 vssd2 vccd2 vccd2 _5969_/B sky130_fd_sc_hd__nor2_1
XANTENNA__6773__A2 _6549_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3895__A _4267_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_90_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4918_ _4919_/A _4919_/B vssd2 vssd2 vccd2 vccd2 _4918_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_47_343 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7706_ _7787_/CLK _7706_/D vssd2 vssd2 vccd2 vccd2 _7706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_62_313 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7637_ _7641_/A vssd2 vssd2 vccd2 vccd2 _7637_/Y sky130_fd_sc_hd__inv_2
X_5898_ _6283_/A _5992_/B _5898_/C vssd2 vssd2 vccd2 vccd2 _5898_/X sky130_fd_sc_hd__and3_1
XFILLER_0_74_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4849_ _4769_/B _4849_/B _4849_/C vssd2 vssd2 vccd2 vccd2 _4997_/A sky130_fd_sc_hd__nand3b_2
XFILLER_0_99_81 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7568_ _7613_/A vssd2 vssd2 vccd2 vccd2 _7568_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
X_6519_ _6519_/A _6519_/B vssd2 vssd2 vccd2 vccd2 _6520_/B sky130_fd_sc_hd__xor2_2
X_7499_ _7561_/A vssd2 vssd2 vccd2 vccd2 _7499_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7486__B1 hold104/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_101_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_100_153 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_100_197 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4892__C _5315_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_85_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_78_490 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4224__B1 _5029_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5972__B1 _6812_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_38_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_93_460 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_81_611 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_108_253 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4527__A1 _4966_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_53_357 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_110_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4527__B2 _4962_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_80_187 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_21_221 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_111_429 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7477__B1 _7483_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_95_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_405 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_66 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_28_88 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_88_221 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_88_265 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6870_ _6871_/B _6871_/A vssd2 vssd2 vccd2 vccd2 _6916_/B sky130_fd_sc_hd__and2b_1
X_5821_ _5821_/A _5821_/B vssd2 vssd2 vccd2 vccd2 _7034_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_48_129 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6803__B _7140_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_57_663 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_8_226 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5752_ _6283_/B _6587_/B vssd2 vssd2 vccd2 vccd2 _5752_/Y sky130_fd_sc_hd__nand2_2
X_4703_ _4704_/B _5142_/C _5076_/D _4898_/A vssd2 vssd2 vccd2 vccd2 _4703_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_44_313 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_29_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_1_0__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_60_97 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_44_357 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5683_ _5735_/B _5682_/X _5679_/X _7879_/Q vssd2 vssd2 vccd2 vccd2 _5944_/B sky130_fd_sc_hd__o2bb2a_4
X_4634_ _4966_/A _4711_/A _5042_/B _4782_/B vssd2 vssd2 vccd2 vccd2 _4635_/B sky130_fd_sc_hd__or4_1
XFILLER_0_8_10 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7422_ _7440_/A _7422_/B vssd2 vssd2 vccd2 vccd2 _7679_/D sky130_fd_sc_hd__and2_1
Xhold612 _7813_/Q vssd2 vssd2 vccd2 vccd2 hold612/X sky130_fd_sc_hd__dlygate4sd3_1
X_4565_ _4565_/A _4565_/B vssd2 vssd2 vccd2 vccd2 _4566_/B sky130_fd_sc_hd__nand2_1
X_7353_ hold153/X _7647_/Q _7383_/S vssd2 vssd2 vccd2 vccd2 _7353_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_43 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold601 hold95/X vssd2 vssd2 vccd2 vccd2 input1/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 hold645/A vssd2 vssd2 vccd2 vccd2 hold645/X sky130_fd_sc_hd__dlygate4sd3_1
X_6304_ _6242_/A _6242_/B _6240_/X vssd2 vssd2 vccd2 vccd2 _6306_/B sky130_fd_sc_hd__a21oi_2
Xhold634 _7820_/Q vssd2 vssd2 vccd2 vccd2 hold634/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 hold623/A vssd2 vssd2 vccd2 vccd2 hold623/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7468__B1 _7483_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold656 _7836_/Q vssd2 vssd2 vccd2 vccd2 hold656/X sky130_fd_sc_hd__dlygate4sd3_1
X_7284_ _7308_/B _7284_/B vssd2 vssd2 vccd2 vccd2 _7310_/C sky130_fd_sc_hd__and2_1
Xhold667 hold667/A vssd2 vssd2 vccd2 vccd2 hold667/X sky130_fd_sc_hd__dlygate4sd3_1
X_4496_ _4704_/B _4896_/A _4711_/A _4782_/B vssd2 vssd2 vccd2 vccd2 _4497_/B sky130_fd_sc_hd__or4_1
Xhold678 _7673_/Q vssd2 vssd2 vccd2 vccd2 hold678/X sky130_fd_sc_hd__dlygate4sd3_1
X_6235_ _6169_/A _6169_/B _6167_/Y vssd2 vssd2 vccd2 vccd2 _6237_/B sky130_fd_sc_hd__a21bo_1
Xhold689 _7665_/Q vssd2 vssd2 vccd2 vccd2 hold689/X sky130_fd_sc_hd__dlygate4sd3_1
X_6166_ _6106_/A _6106_/B _6106_/C vssd2 vssd2 vccd2 vccd2 _6168_/B sky130_fd_sc_hd__a21boi_2
XTAP_961 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6266__A _6855_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5117_ _5118_/A _5118_/B vssd2 vssd2 vccd2 vccd2 _5117_/Y sky130_fd_sc_hd__nor2_1
XTAP_994 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _7847_/Q _6510_/B _6670_/B _7846_/Q vssd2 vssd2 vccd2 vccd2 _6097_/X sky130_fd_sc_hd__a22o_1
X_5048_ _5048_/A _5048_/B vssd2 vssd2 vccd2 vccd2 _5051_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__6416__D _6973_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_79_221 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6713__B _7181_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7097__A _7143_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6999_ _6999_/A _6999_/B vssd2 vssd2 vccd2 vccd2 _7001_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_75_482 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_75_460 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_47_173 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_90_441 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_63_655 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_35_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_105_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_90_463 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_62_176 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_7_270 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_62_187 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7459__B1 _7485_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_31_585 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_101_462 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__6434__A1 _6253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_105_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_58_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_14_24 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_85_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_38_151 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_38_162 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_109_584 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_38_184 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_14_508 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_26_379 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_30_78 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_30_89 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4350_ _4350_/A _4350_/B vssd2 vssd2 vccd2 vccd2 _4351_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_111_237 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_1_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4281_ _5042_/A _5029_/A vssd2 vssd2 vccd2 vccd2 _4283_/A sky130_fd_sc_hd__or2_2
XFILLER_0_39_54 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_65 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_257 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6020_ _7850_/Q _5791_/X _6014_/X _6016_/X _6018_/X vssd2 vssd2 vccd2 vccd2 _6020_/X
+ sky130_fd_sc_hd__a2111o_2
XTAP_268 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_530 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_55_97 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6922_ _6922_/A _6922_/B vssd2 vssd2 vccd2 vccd2 _6925_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_89_596 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_71_30 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6853_ _6854_/A _6854_/B vssd2 vssd2 vccd2 vccd2 _6853_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_49_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_49_438 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_64_408 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_9_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5804_ _7847_/Q _6075_/C _6075_/D _7843_/Q _5659_/B vssd2 vssd2 vccd2 vccd2 _5804_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_91_205 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6784_ _6784_/A _6784_/B vssd2 vssd2 vccd2 vccd2 _6795_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__4334__A _4962_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3996_ _4328_/A _3996_/B _4268_/D _4002_/B vssd2 vssd2 vccd2 vccd2 _3996_/X sky130_fd_sc_hd__and4_1
XANTENNA__7348__C _7385_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_29_173 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_91_249 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_72_441 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_72_430 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_57_493 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_45_633 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_44_132 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5735_ _7871_/Q _5735_/B vssd2 vssd2 vccd2 vccd2 _5736_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_95_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_60_603 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5666_ _6282_/A _5878_/B _5836_/B _5665_/Y vssd2 vssd2 vccd2 vccd2 _5666_/X sky130_fd_sc_hd__a22o_1
X_4617_ _4617_/A _4617_/B vssd2 vssd2 vccd2 vccd2 _4618_/B sky130_fd_sc_hd__xnor2_2
X_7405_ _7452_/A _7405_/B vssd2 vssd2 vccd2 vccd2 _7405_/X sky130_fd_sc_hd__and2_1
Xhold420 la_data_in[41] vssd2 vssd2 vccd2 vccd2 hold1/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5165__A _5220_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5597_ _7867_/Q _5598_/B vssd2 vssd2 vccd2 vccd2 _5659_/B sky130_fd_sc_hd__xor2_4
XANTENNA__6361__B1 _6281_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7336_ _7336_/A _7336_/B vssd2 vssd2 vccd2 vccd2 _7838_/D sky130_fd_sc_hd__and2_1
Xhold453 hold25/X vssd2 vssd2 vccd2 vccd2 input41/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 input33/X vssd2 vssd2 vccd2 vccd2 hold10/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 hold6/X vssd2 vssd2 vccd2 vccd2 _7881_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4548_ _4420_/A _4420_/B _4480_/C _4422_/A vssd2 vssd2 vccd2 vccd2 _4551_/B sky130_fd_sc_hd__a211o_1
X_7267_ _7267_/A _7267_/B vssd2 vssd2 vccd2 vccd2 _7268_/B sky130_fd_sc_hd__and2_1
Xhold464 la_data_in[40] vssd2 vssd2 vccd2 vccd2 hold23/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 input6/X vssd2 vssd2 vccd2 vccd2 hold22/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 hold42/X vssd2 vssd2 vccd2 vccd2 _7857_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4479_ _4479_/A _4479_/B vssd2 vssd2 vccd2 vccd2 _4480_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__5315__D _5468_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6218_ _6668_/A _7047_/A vssd2 vssd2 vccd2 vccd2 _6229_/A sky130_fd_sc_hd__nand2_1
Xhold497 hold51/X vssd2 vssd2 vccd2 vccd2 input9/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7380__A _7452_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5467__A2 _5528_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7198_ _7199_/B _7199_/C _7199_/A vssd2 vssd2 vccd2 vccd2 _7242_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_99_305 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6149_ _6149_/A _6149_/B vssd2 vssd2 vccd2 vccd2 _6169_/A sky130_fd_sc_hd__xor2_2
XTAP_791 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_349 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_95_544 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_82_205 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_35_121 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7555__A _7563_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_50_124 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4898__B _5528_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_23_327 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_35_187 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_50_146 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6104__B1 _7047_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_31_382 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_31_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_101_281 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_92_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_46_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3850_ _7793_/Q _3851_/B vssd2 vssd2 vccd2 vccd2 _4083_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_39_471 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_41_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_54_474 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_14_305 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5520_ _5488_/A _5485_/Y _5486_/X vssd2 vssd2 vccd2 vccd2 _5522_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_41_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_112_513 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5451_ _5451_/A _5451_/B vssd2 vssd2 vccd2 vccd2 _5453_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_112_557 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4402_ _4402_/A _4402_/B vssd2 vssd2 vccd2 vccd2 _4404_/B sky130_fd_sc_hd__xnor2_4
X_5382_ _5382_/A _5382_/B vssd2 vssd2 vccd2 vccd2 _5385_/A sky130_fd_sc_hd__xnor2_4
X_7121_ _7121_/A _7121_/B vssd2 vssd2 vccd2 vccd2 _7123_/B sky130_fd_sc_hd__xnor2_1
X_4333_ _4810_/A _5099_/A vssd2 vssd2 vccd2 vccd2 _4338_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_10_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_22_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xfanout207 _4129_/Y vssd2 vssd2 vccd2 vccd2 _5029_/A sky130_fd_sc_hd__clkbuf_8
X_7052_ _7052_/A _7052_/B vssd2 vssd2 vccd2 vccd2 _7054_/A sky130_fd_sc_hd__xor2_2
Xfanout229 _7485_/B1 vssd2 vssd2 vccd2 vccd2 _7483_/B1 sky130_fd_sc_hd__buf_4
XANTENNA__7404__S _7418_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4264_ _4262_/Y _4263_/X _4745_/A vssd2 vssd2 vccd2 vccd2 _4264_/Y sky130_fd_sc_hd__a21oi_1
Xfanout218 _4628_/X vssd2 vssd2 vccd2 vccd2 _5498_/A sky130_fd_sc_hd__buf_4
X_6003_ _6003_/A _6003_/B _6003_/C vssd2 vssd2 vccd2 vccd2 _6003_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_66_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4195_ _4196_/A _4195_/B vssd2 vssd2 vccd2 vccd2 _7731_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__7071__A1 _6989_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6905_ _7025_/C vssd2 vssd2 vccd2 vccd2 _6908_/A sky130_fd_sc_hd__inv_2
XFILLER_0_89_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_82_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1209 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_10_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA_fanout266_A _7806_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3887__B _4267_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7885_ _7886_/CLK _7885_/D _7644_/Y vssd2 vssd2 vccd2 vccd2 _7885_/Q sky130_fd_sc_hd__dfrtp_4
X_6836_ _6839_/A _6839_/B vssd2 vssd2 vccd2 vccd2 _6836_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_49_268 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_37_408 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6767_ _6767_/A _6767_/B _6767_/C vssd2 vssd2 vccd2 vccd2 _6768_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_9_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4999__A _5133_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_17_110 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_107_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5718_ _7873_/Q _7872_/Q _7871_/Q _7874_/Q _5735_/B vssd2 vssd2 vccd2 vccd2 _5731_/B
+ sky130_fd_sc_hd__o41a_2
X_3979_ _3945_/Y _3975_/X _3976_/X _3978_/X vssd2 vssd2 vccd2 vccd2 _3979_/X sky130_fd_sc_hd__a31o_1
X_6698_ _6637_/A _6637_/B _6635_/B vssd2 vssd2 vccd2 vccd2 _6700_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_72_260 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_17_198 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_103_524 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_103_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5649_ _5661_/B _5836_/B _5649_/C vssd2 vssd2 vccd2 vccd2 _5807_/C sky130_fd_sc_hd__and3_1
Xhold261 hold614/X vssd2 vssd2 vccd2 vccd2 hold615/A sky130_fd_sc_hd__dlygate4sd3_1
X_7319_ _7319_/A _7319_/B _7319_/C vssd2 vssd2 vccd2 vccd2 _7320_/B sky130_fd_sc_hd__nand3_1
Xhold250 _7455_/X vssd2 vssd2 vccd2 vccd2 _7695_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 hold272/A vssd2 vssd2 vccd2 vccd2 la_data_out[30] sky130_fd_sc_hd__buf_12
Xhold294 hold294/A vssd2 vssd2 vccd2 vccd2 la_data_out[20] sky130_fd_sc_hd__buf_12
Xhold283 hold636/X vssd2 vssd2 vccd2 vccd2 hold637/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_113 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_68_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_68_511 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_68_555 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_83_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_68_577 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_83_558 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6573__B1 _6150_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_249 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_102_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_51_466 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_51_433 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6629__A _6670_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xinput7 input7/A vssd2 vssd2 vccd2 vccd2 input7/X sky130_fd_sc_hd__buf_1
XANTENNA__5851__A2 _6281_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_36_22 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4951_ _4951_/A _4951_/B vssd2 vssd2 vccd2 vccd2 _4982_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_86_352 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_74_525 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4882_ _4882_/A _5164_/B _4883_/A vssd2 vssd2 vccd2 vccd2 _4882_/X sky130_fd_sc_hd__or3_1
X_7670_ _7782_/CLK _7670_/D vssd2 vssd2 vccd2 vccd2 _7670_/Q sky130_fd_sc_hd__dfxtp_1
X_3902_ _4148_/C _4148_/D _3902_/C _4010_/D vssd2 vssd2 vccd2 vccd2 _3902_/Y sky130_fd_sc_hd__nor4_1
X_6621_ _6769_/A _6769_/B _7034_/A vssd2 vssd2 vccd2 vccd2 _6696_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_558 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_46_249 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_46_227 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3833_ _7799_/Q _3822_/A _3822_/B _3888_/B vssd2 vssd2 vccd2 vccd2 _3835_/B sky130_fd_sc_hd__o31a_2
XANTENNA__5367__A1 _5366_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_61_219 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_54_271 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6552_ _5945_/X _5947_/X _7143_/B _5755_/C vssd2 vssd2 vccd2 vccd2 _6556_/A sky130_fd_sc_hd__o211a_2
X_6483_ _6483_/A _6483_/B vssd2 vssd2 vccd2 vccd2 _6486_/A sky130_fd_sc_hd__or2_1
XANTENNA__4590__A2 _5042_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_15_647 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5503_ _5503_/A _5503_/B vssd2 vssd2 vccd2 vccd2 _5506_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_321 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_42_499 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_42_488 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5434_ _5480_/B _5436_/B vssd2 vssd2 vccd2 vccd2 _5437_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_112_365 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_100_549 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7104_ _7104_/A _7104_/B vssd2 vssd2 vccd2 vccd2 _7106_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5365_ _5365_/A _5365_/B vssd2 vssd2 vccd2 vccd2 _5366_/C sky130_fd_sc_hd__xor2_1
X_5296_ _5294_/X _5296_/B vssd2 vssd2 vccd2 vccd2 _5297_/B sky130_fd_sc_hd__nand2b_1
X_4316_ _7768_/Q _4707_/A _4063_/X _4162_/A vssd2 vssd2 vccd2 vccd2 _4316_/X sky130_fd_sc_hd__a22o_1
X_7035_ _7131_/A _7035_/B vssd2 vssd2 vccd2 vccd2 _7827_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__7292__A1 _7253_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7292__B2 _7253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4247_ _4303_/A _4247_/B vssd2 vssd2 vccd2 vccd2 _4305_/B sky130_fd_sc_hd__xnor2_1
X_4178_ _4178_/A _4178_/B vssd2 vssd2 vccd2 vccd2 _4180_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__7044__B2 _7094_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7044__A1 _7197_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6705__C _7253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1028 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_216 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7868_ _7870_/CLK _7868_/D _7627_/Y vssd2 vssd2 vccd2 vccd2 _7868_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_92_333 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6819_ _6819_/A _6819_/B vssd2 vssd2 vccd2 vccd2 _6820_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_151 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_80_506 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7799_ _7802_/CLK _7799_/D _7558_/Y vssd2 vssd2 vccd2 vccd2 _7799_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5618__A _7844_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_107_137 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_80_528 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_45_260 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4522__A _7772_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_45_293 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_60_274 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_60_263 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_33_499 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_87_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XTAP_1551 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1584 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_193 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_91 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_22_24 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_28_249 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_80 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_377 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_22_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5528__A _5528_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_83_388 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_71_528 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_36_282 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_24_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5150_ _5276_/A _5414_/A vssd2 vssd2 vccd2 vccd2 _5154_/B sky130_fd_sc_hd__nor2_1
X_5081_ _5210_/A _5210_/B _5081_/C _5468_/A vssd2 vssd2 vccd2 vccd2 _5082_/B sky130_fd_sc_hd__or4_1
XFILLER_0_47_54 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4101_ _4101_/A vssd2 vssd2 vccd2 vccd2 _4101_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_87 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4032_ _7763_/Q _4033_/C _4032_/C vssd2 vssd2 vccd2 vccd2 _4032_/X sky130_fd_sc_hd__and3_1
XANTENNA__6094__A _6158_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6785__B1 _7143_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5983_ _5975_/X _5977_/X _5980_/X _5981_/X _5811_/C vssd2 vssd2 vccd2 vccd2 _5984_/B
+ sky130_fd_sc_hd__o41ai_4
X_4934_ _5042_/B _5404_/A vssd2 vssd2 vccd2 vccd2 _4935_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_63_86 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_59_374 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7722_ _7723_/CLK _7722_/D vssd2 vssd2 vccd2 vccd2 _7722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_333 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_59_385 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7329__A2 _7197_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_19_wb_clk_i clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7779_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_216 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4865_ _5210_/B _4965_/B _5222_/A _5210_/A vssd2 vssd2 vccd2 vccd2 _4865_/X sky130_fd_sc_hd__o22a_1
X_7653_ _7779_/CLK _7653_/D vssd2 vssd2 vccd2 vccd2 _7653_/Q sky130_fd_sc_hd__dfxtp_1
X_7584_ _7590_/A vssd2 vssd2 vccd2 vccd2 _7584_/Y sky130_fd_sc_hd__inv_2
X_6604_ _6604_/A _6604_/B vssd2 vssd2 vccd2 vccd2 _6607_/A sky130_fd_sc_hd__xnor2_2
X_4796_ _5029_/A _5406_/A vssd2 vssd2 vccd2 vccd2 _4799_/A sky130_fd_sc_hd__or2_1
XANTENNA__4342__A _5029_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_7_644 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA_fanout229_A _7485_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3816_ _7803_/Q _3822_/A _3822_/B _3822_/C _3888_/B vssd2 vssd2 vccd2 vccd2 _3818_/B
+ sky130_fd_sc_hd__o41a_4
XANTENNA__4012__B2 _7764_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6535_ _6536_/B _6536_/A vssd2 vssd2 vccd2 vccd2 _6613_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_103_81 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4563__A2 _4711_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_113_630 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_42_241 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6466_ _6466_/A _6466_/B vssd2 vssd2 vccd2 vccd2 _6467_/B sky130_fd_sc_hd__or2_1
XANTENNA__4996__B _4996_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_30_425 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_88_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xoutput130 hold611/X vssd2 vssd2 vccd2 vccd2 hold258/A sky130_fd_sc_hd__buf_6
X_6397_ _6397_/A _7313_/A vssd2 vssd2 vccd2 vccd2 _6397_/Y sky130_fd_sc_hd__nand2_1
Xoutput141 _7711_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[16] sky130_fd_sc_hd__buf_12
Xoutput152 _7721_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[26] sky130_fd_sc_hd__buf_12
XFILLER_0_2_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5417_ _5417_/A _5417_/B vssd2 vssd2 vccd2 vccd2 _5418_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_112_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5348_ _5349_/A _5349_/B vssd2 vssd2 vccd2 vccd2 _5395_/B sky130_fd_sc_hd__or2_1
Xoutput163 _7702_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[7] sky130_fd_sc_hd__buf_12
XANTENNA__7265__B2 _7291_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7018_ _7019_/A _7019_/B vssd2 vssd2 vccd2 vccd2 _7081_/B sky130_fd_sc_hd__nor2_1
X_5279_ _5279_/A _5279_/B vssd2 vssd2 vccd2 vccd2 _5281_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_311 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_92_141 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_65_388 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_104_641 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_61_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7563__A _7563_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5083__A _5366_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_609 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7008__A1 _6939_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_88_425 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_17_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_88_469 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6642__A _6855_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_8_408 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1392 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5990__A1 _7847_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4650_ _4729_/A _4965_/B _5030_/B vssd2 vssd2 vccd2 vccd2 _4651_/B sky130_fd_sc_hd__or3b_2
XANTENNA__7176__C _7291_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_56_399 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__4162__A _4162_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_114_405 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_71_358 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xinput10 input10/A vssd2 vssd2 vccd2 vccd2 input10/X sky130_fd_sc_hd__clkbuf_1
Xinput21 input21/A vssd2 vssd2 vccd2 vccd2 input21/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_449 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6320_ _6387_/B _6320_/B vssd2 vssd2 vccd2 vccd2 _6390_/B sky130_fd_sc_hd__nand2_1
X_4581_ _4581_/A _4581_/B vssd2 vssd2 vccd2 vccd2 _4583_/B sky130_fd_sc_hd__xnor2_2
Xinput32 input32/A vssd2 vssd2 vccd2 vccd2 input32/X sky130_fd_sc_hd__clkbuf_1
Xinput43 input43/A vssd2 vssd2 vccd2 vccd2 input43/X sky130_fd_sc_hd__clkbuf_1
Xinput54 wbs_adr_i[13] vssd2 vssd2 vccd2 vccd2 _7343_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xinput98 input98/A vssd2 vssd2 vccd2 vccd2 input98/X sky130_fd_sc_hd__clkbuf_1
Xinput87 input87/A vssd2 vssd2 vccd2 vccd2 input87/X sky130_fd_sc_hd__clkbuf_1
Xinput65 wbs_adr_i[23] vssd2 vssd2 vccd2 vccd2 _7340_/C sky130_fd_sc_hd__clkbuf_1
Xinput76 wbs_adr_i[4] vssd2 vssd2 vccd2 vccd2 _7342_/B sky130_fd_sc_hd__clkbuf_1
X_6251_ _6402_/A _7143_/A vssd2 vssd2 vccd2 vccd2 _6259_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6089__A _6812_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6182_ _6182_/A _6182_/B vssd2 vssd2 vccd2 vccd2 _6185_/A sky130_fd_sc_hd__xnor2_2
X_5202_ _5168_/A _5431_/B _5301_/A _5201_/X vssd2 vssd2 vccd2 vccd2 _5240_/A sky130_fd_sc_hd__o22ai_4
XFILLER_0_58_42 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5133_ _5133_/A _5133_/B _5133_/C _5133_/D vssd2 vssd2 vccd2 vccd2 _5357_/A sky130_fd_sc_hd__nand4_2
XFILLER_0_20_491 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7412__S _7418_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5721__A _5992_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5064_ _5064_/A _5064_/B vssd2 vssd2 vccd2 vccd2 _5067_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_74_41 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6470__A2 _7222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_74_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_74_63 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4015_ _7766_/Q _4075_/B _4200_/B _7768_/Q _3996_/X vssd2 vssd2 vccd2 vccd2 _4015_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_0_79_436 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA_fanout179_A _6642_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_480 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5966_ _6064_/A _5966_/B vssd2 vssd2 vccd2 vccd2 _5968_/A sky130_fd_sc_hd__nand2_1
X_4917_ _4834_/A _4834_/B _4832_/Y vssd2 vssd2 vccd2 vccd2 _4919_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_74_141 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5981__A1 _6157_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5981__B2 _7847_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7705_ _7802_/CLK _7705_/D vssd2 vssd2 vccd2 vccd2 _7705_/Q sky130_fd_sc_hd__dfxtp_1
X_5897_ _7843_/Q _6588_/B _5751_/Y _7844_/Q vssd2 vssd2 vccd2 vccd2 _5897_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_47_366 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__5168__A _5168_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4848_ _4849_/B _4848_/B vssd2 vssd2 vccd2 vccd2 _7741_/D sky130_fd_sc_hd__xor2_2
X_7636_ _7641_/A vssd2 vssd2 vccd2 vccd2 _7636_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_430 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_105_405 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_105_449 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4779_ _4779_/A _5550_/A vssd2 vssd2 vccd2 vccd2 _4780_/B sky130_fd_sc_hd__nor2_2
X_7567_ _7613_/A vssd2 vssd2 vccd2 vccd2 _7567_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_572 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_43_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_99_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6518_ _6519_/A _6519_/B vssd2 vssd2 vccd2 vccd2 _6518_/X sky130_fd_sc_hd__and2_1
XFILLER_0_70_380 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4800__A _5030_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7498_ _7524_/A vssd2 vssd2 vccd2 vccd2 _7498_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_274 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6449_ _6449_/A _6449_/B vssd2 vssd2 vccd2 vccd2 _6450_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_100_121 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5497__B1 _5498_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_30_288 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_100_165 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_11_491 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_11_480 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_30_299 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_85_439 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5972__A1 _5778_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_108_221 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_93_472 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5078__A _5168_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_26_528 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_38_388 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_108_265 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_53_369 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6921__B1 _7294_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_41_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_110_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_406 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_233 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_88_277 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__3996__A _4328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5820_ _7886_/Q _5821_/B vssd2 vssd2 vccd2 vccd2 _5820_/X sky130_fd_sc_hd__xor2_1
XANTENNA__4215__A1 _4268_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_91_409 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_56_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5751_ _6100_/D _6510_/B vssd2 vssd2 vccd2 vccd2 _5751_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_84_472 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4702_ _4655_/A _4653_/Y _4652_/Y vssd2 vssd2 vccd2 vccd2 _4720_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_44_347 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5682_ _5694_/A _5694_/B _5694_/C _7879_/Q vssd2 vssd2 vccd2 vccd2 _5682_/X sky130_fd_sc_hd__o31a_1
X_7421_ hold153/X _7791_/D _7451_/S vssd2 vssd2 vccd2 vccd2 _7421_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6912__B1 _7034_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4633_ _4711_/A _5042_/B _4782_/B _4966_/A vssd2 vssd2 vccd2 vccd2 _4633_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_71_155 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_44_369 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5716__A _7847_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4564_ _4896_/A _4966_/A _4711_/A _4782_/B vssd2 vssd2 vccd2 vccd2 _4565_/B sky130_fd_sc_hd__or4_1
Xhold602 input1/X vssd2 vssd2 vccd2 vccd2 hold96/A sky130_fd_sc_hd__dlygate4sd3_1
X_7352_ _7454_/A _7420_/A vssd2 vssd2 vccd2 vccd2 _7352_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_520 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold624 _7828_/Q vssd2 vssd2 vccd2 vccd2 hold624/X sky130_fd_sc_hd__dlygate4sd3_1
X_6303_ _6303_/A _6303_/B vssd2 vssd2 vccd2 vccd2 _6306_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7283_ _7283_/A _7283_/B _7283_/C vssd2 vssd2 vccd2 vccd2 _7284_/B sky130_fd_sc_hd__nand3_1
Xhold635 hold635/A vssd2 vssd2 vccd2 vccd2 hold635/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 hold613/A vssd2 vssd2 vccd2 vccd2 hold613/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold657 hold657/A vssd2 vssd2 vccd2 vccd2 hold657/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 _7835_/Q vssd2 vssd2 vccd2 vccd2 hold668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 _7822_/Q vssd2 vssd2 vccd2 vccd2 hold646/X sky130_fd_sc_hd__dlygate4sd3_1
X_6234_ _6234_/A _6234_/B vssd2 vssd2 vccd2 vccd2 _6237_/A sky130_fd_sc_hd__xnor2_2
X_4495_ _4896_/A _4711_/A _4782_/B _4704_/B vssd2 vssd2 vccd2 vccd2 _4497_/A sky130_fd_sc_hd__o22ai_1
XFILLER_0_12_277 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold679 _7651_/Q vssd2 vssd2 vccd2 vccd2 hold679/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_474 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_85_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6165_ _6165_/A _6165_/B vssd2 vssd2 vccd2 vccd2 _6168_/A sky130_fd_sc_hd__xnor2_2
XTAP_951 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5451__A _5451_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_40_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6266__B _6973_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5116_ _5056_/A _5056_/B _5054_/X vssd2 vssd2 vccd2 vccd2 _5118_/B sky130_fd_sc_hd__a21oi_2
XTAP_995 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _6094_/Y _6095_/X _6283_/B _6510_/B vssd2 vssd2 vccd2 vccd2 _6096_/Y sky130_fd_sc_hd__a211oi_1
X_5047_ _5047_/A _5047_/B vssd2 vssd2 vccd2 vccd2 _5048_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_67_406 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7378__A _7452_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6282__A _6282_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6998_ _6986_/A _7181_/A _6946_/A _6943_/Y vssd2 vssd2 vccd2 vccd2 _6999_/B sky130_fd_sc_hd__o31ai_2
XANTENNA__5954__A1 _6402_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7097__B _7143_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5949_ _5945_/X _5947_/X _5755_/C vssd2 vssd2 vccd2 vccd2 _6705_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__5403__B1 _5498_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_47_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_303 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7156__B1 _7037_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_62_122 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_90_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_62_166 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7619_ _7645_/A vssd2 vssd2 vccd2 vccd2 _7619_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_35_369 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_50_328 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_105_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6131__B2 _7850_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6131__A1 _6670_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_98_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_105_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_98_597 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_85_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5945__A1 _6283_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5945__B2 _6158_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_38_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_109_574 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_54_645 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_30_13 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_81_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7454__C _7454_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_22_520 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_41_328 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_111_205 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5255__B _5357_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_22_542 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_111_249 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_39_22 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_4280_ _4729_/A _4863_/A _5030_/B vssd2 vssd2 vccd2 vccd2 _4285_/A sky130_fd_sc_hd__or3b_2
XFILLER_0_39_44 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XTAP_236 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_87 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_55_54 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5633__B1 _5645_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6921_ _6020_/X _6021_/X _7294_/C _5811_/B vssd2 vssd2 vccd2 vccd2 _6922_/B sky130_fd_sc_hd__o211a_1
X_6852_ _6039_/X _6040_/X _7222_/A _5992_/B vssd2 vssd2 vccd2 vccd2 _6854_/B sky130_fd_sc_hd__o211a_1
XFILLER_0_71_42 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_9_525 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5803_ _6253_/B _6018_/D _5835_/D _5803_/D vssd2 vssd2 vccd2 vccd2 _5803_/X sky130_fd_sc_hd__and4_1
XFILLER_0_91_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6783_ _6783_/A _7255_/B vssd2 vssd2 vccd2 vccd2 _6784_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4334__B _4966_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3995_ _3996_/B _4268_/D _4002_/B vssd2 vssd2 vccd2 vccd2 _3995_/X sky130_fd_sc_hd__and3_1
XANTENNA__3876__D _4267_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5734_ _7873_/Q _5734_/B vssd2 vssd2 vccd2 vccd2 _5734_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_72_464 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_44_166 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_44_155 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5665_ _6587_/A _5665_/B _5812_/C vssd2 vssd2 vccd2 vccd2 _5665_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_88_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4616_ _4617_/A _4617_/B vssd2 vssd2 vccd2 vccd2 _4685_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_44_188 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7404_ hold121/X _7671_/Q _7418_/S vssd2 vssd2 vccd2 vccd2 _7404_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_520 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_32_317 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_111_81 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7335_ _7335_/A _7335_/B _7334_/X vssd2 vssd2 vccd2 vccd2 _7336_/B sky130_fd_sc_hd__or3b_4
X_5596_ _7868_/Q _5598_/B vssd2 vssd2 vccd2 vccd2 _5599_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__5165__B _5406_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_25_391 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold410 _7886_/Q vssd2 vssd2 vccd2 vccd2 _5821_/A sky130_fd_sc_hd__clkbuf_2
Xhold454 input41/X vssd2 vssd2 vccd2 vccd2 hold26/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 hold1/X vssd2 vssd2 vccd2 vccd2 input36/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 la_data_in[37] vssd2 vssd2 vccd2 vccd2 hold33/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 hold10/X vssd2 vssd2 vccd2 vccd2 _7846_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4547_ _4547_/A _4547_/B vssd2 vssd2 vccd2 vccd2 _4551_/A sky130_fd_sc_hd__xnor2_2
Xmax_cap184 _6873_/A vssd2 vssd2 vccd2 vccd2 _6581_/A sky130_fd_sc_hd__buf_2
X_7266_ _7267_/A _7267_/B vssd2 vssd2 vccd2 vccd2 _7300_/A sky130_fd_sc_hd__nor2_1
Xhold465 hold23/X vssd2 vssd2 vccd2 vccd2 input35/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 hold22/X vssd2 vssd2 vccd2 vccd2 _7885_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 la_data_in[20] vssd2 vssd2 vccd2 vccd2 hold13/A sky130_fd_sc_hd__dlygate4sd3_1
X_4478_ _4478_/A _4478_/B vssd2 vssd2 vccd2 vccd2 _4479_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6217_ _6217_/A _6217_/B vssd2 vssd2 vccd2 vccd2 _6234_/A sky130_fd_sc_hd__xor2_2
X_7197_ _7197_/A _7197_/B vssd2 vssd2 vccd2 vccd2 _7199_/C sky130_fd_sc_hd__nand2_1
Xhold498 input9/X vssd2 vssd2 vccd2 vccd2 hold52/A sky130_fd_sc_hd__dlygate4sd3_1
X_6148_ _6148_/A _6148_/B vssd2 vssd2 vccd2 vccd2 _6149_/B sky130_fd_sc_hd__nand2_1
XTAP_770 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_317 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4509__B _5042_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_792 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _6073_/Y _6920_/A2 _5664_/C vssd2 vssd2 vccd2 vccd2 _6571_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_95_523 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4525__A _5315_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_67_247 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__5927__B2 _7846_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5927__A1 _6158_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3938__B1 _4050_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_36_645 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_106_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_63_464 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_63_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_144 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_177 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_35_199 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_50_136 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7571__A _7613_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_101_293 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6634__B _6634_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_25_24 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_26_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_39_483 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_54_442 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_41_78 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_109_393 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5450_ _4996_/B _5249_/X _5448_/Y _5449_/Y vssd2 vssd2 vccd2 vccd2 _5451_/B sky130_fd_sc_hd__a31oi_4
XFILLER_0_112_525 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4401_ _4401_/A _4401_/B vssd2 vssd2 vccd2 vccd2 _4402_/B sky130_fd_sc_hd__xnor2_4
X_5381_ _5381_/A _5381_/B vssd2 vssd2 vccd2 vccd2 _5382_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7120_ _7166_/B _7120_/B _7121_/B vssd2 vssd2 vccd2 vccd2 _7169_/A sky130_fd_sc_hd__or3_1
X_4332_ _4327_/X _4331_/X _4267_/D vssd2 vssd2 vccd2 vccd2 _5207_/A sky130_fd_sc_hd__o21ai_4
Xfanout219 _4628_/X vssd2 vssd2 vccd2 vccd2 _5076_/D sky130_fd_sc_hd__clkbuf_4
X_7051_ _7051_/A _7224_/A _7052_/B vssd2 vssd2 vccd2 vccd2 _7051_/X sky130_fd_sc_hd__or3_1
Xfanout208 _4704_/B vssd2 vssd2 vccd2 vccd2 _5042_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_556 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4263_ _3813_/A _3813_/B _4454_/B _3886_/C _4490_/A vssd2 vssd2 vccd2 vccd2 _4263_/X
+ sky130_fd_sc_hd__a2111o_1
X_6002_ _6001_/A _6001_/B _6001_/C vssd2 vssd2 vccd2 vccd2 _6003_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_10_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4657__A1 _4268_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4194_ _5548_/A _4196_/B vssd2 vssd2 vccd2 vccd2 _4195_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_96_309 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_82_41 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__7071__A2 _7291_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6904_ _6904_/A _6904_/B vssd2 vssd2 vccd2 vccd2 _7025_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_82_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_77_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_49_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7884_ _7886_/CLK _7884_/D _7643_/Y vssd2 vssd2 vccd2 vccd2 _7884_/Q sky130_fd_sc_hd__dfrtp_4
X_6835_ _6839_/A _6839_/B vssd2 vssd2 vccd2 vccd2 _6838_/A sky130_fd_sc_hd__and2_1
X_6766_ _6461_/A _6461_/B _6765_/A _6615_/Y _6765_/C vssd2 vssd2 vccd2 vccd2 _6767_/C
+ sky130_fd_sc_hd__a2111o_2
XFILLER_0_92_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_9_377 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3978_ _7765_/Q _4814_/B _4315_/B _4022_/B _3977_/X vssd2 vssd2 vccd2 vccd2 _3978_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_72_250 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5717_ _6157_/A _5992_/B _5712_/X _5716_/X vssd2 vssd2 vccd2 vccd2 _5717_/X sky130_fd_sc_hd__a31o_1
X_6697_ _6648_/A _6648_/B _6651_/A vssd2 vssd2 vccd2 vccd2 _6700_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_272 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_60_412 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_5_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5648_ _5665_/B _5648_/B vssd2 vssd2 vccd2 vccd2 _5649_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_32_125 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_536 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7391__A _7436_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5579_ _7863_/Q _7864_/Q vssd2 vssd2 vccd2 vccd2 _5579_/X sky130_fd_sc_hd__or2_1
Xhold262 hold262/A vssd2 vssd2 vccd2 vccd2 la_data_out[1] sky130_fd_sc_hd__buf_12
X_7318_ _7319_/A _7319_/B _7319_/C vssd2 vssd2 vccd2 vccd2 _7334_/A sky130_fd_sc_hd__a21o_1
Xhold251 _7728_/Q vssd2 vssd2 vccd2 vccd2 hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 _7460_/X vssd2 vssd2 vccd2 vccd2 _7700_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 hold624/X vssd2 vssd2 vccd2 vccd2 hold625/A sky130_fd_sc_hd__dlygate4sd3_1
X_7249_ _7279_/B _7249_/B vssd2 vssd2 vccd2 vccd2 _7310_/B sky130_fd_sc_hd__xor2_2
Xhold284 hold284/A vssd2 vssd2 vccd2 vccd2 la_data_out[18] sky130_fd_sc_hd__buf_12
Xhold295 hold648/X vssd2 vssd2 vccd2 vccd2 hold649/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_125 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_99_169 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5073__A1 _5042_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_68_523 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_68_589 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7566__A _7613_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_36_453 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_11_48 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_51_456 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_51_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_23_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xinput8 input8/A vssd2 vssd2 vccd2 vccd2 input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_512 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4950_ _4950_/A _4950_/B vssd2 vssd2 vccd2 vccd2 _4951_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_59_545 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_52_33 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_74_504 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4881_ wire212/X _4881_/A2 _5498_/D vssd2 vssd2 vccd2 vccd2 _4883_/B sky130_fd_sc_hd__a21oi_1
X_3901_ _4148_/B _3901_/B vssd2 vssd2 vccd2 vccd2 _4010_/D sky130_fd_sc_hd__nand2_1
X_6620_ _6769_/A _6620_/B vssd2 vssd2 vccd2 vccd2 _7821_/D sky130_fd_sc_hd__xnor2_1
X_3832_ _3822_/A _3822_/B _3888_/B vssd2 vssd2 vccd2 vccd2 _3838_/B sky130_fd_sc_hd__o21a_2
XANTENNA__5367__A2 _5498_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6551_ _6551_/A _6551_/B vssd2 vssd2 vccd2 vccd2 _6563_/A sky130_fd_sc_hd__xnor2_1
X_5502_ _5503_/A _5503_/B vssd2 vssd2 vccd2 vccd2 _5539_/A sky130_fd_sc_hd__nor2_1
X_6482_ _6481_/A _6481_/B _6481_/C vssd2 vssd2 vccd2 vccd2 _6483_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_112_333 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5433_ _5433_/A _5433_/B _5433_/C vssd2 vssd2 vccd2 vccd2 _5436_/B sky130_fd_sc_hd__nor3_1
XANTENNA__5724__A _6152_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5364_ _5414_/A _5550_/A vssd2 vssd2 vccd2 vccd2 _5365_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_112_377 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_100_528 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7103_ _7103_/A _7103_/B vssd2 vssd2 vccd2 vccd2 _7104_/B sky130_fd_sc_hd__xor2_1
X_4315_ _4809_/A _4315_/B _4315_/C _4427_/A vssd2 vssd2 vccd2 vccd2 _4315_/X sky130_fd_sc_hd__and4_1
X_5295_ _5295_/A _5295_/B _5293_/Y vssd2 vssd2 vccd2 vccd2 _5296_/B sky130_fd_sc_hd__or3b_1
XANTENNA__5827__B1 _7846_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7034_ _7034_/A _7326_/A vssd2 vssd2 vccd2 vccd2 _7035_/B sky130_fd_sc_hd__nor2_1
X_4246_ _4303_/A _4247_/B vssd2 vssd2 vccd2 vccd2 _4304_/A sky130_fd_sc_hd__or2_1
XFILLER_0_93_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__6555__A _6556_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4177_ _4177_/A _4177_/B vssd2 vssd2 vccd2 vccd2 _4178_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__7044__A2 _7222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6705__D _7253_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_96_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1029 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4075__A _7767_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_92_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7867_ _7870_/CLK _7867_/D _7626_/Y vssd2 vssd2 vccd2 vccd2 _7867_/Q sky130_fd_sc_hd__dfrtp_4
X_6818_ _6819_/A _6819_/B vssd2 vssd2 vccd2 vccd2 _6818_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_107_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_92_345 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7798_ _7798_/CLK _7798_/D _7557_/Y vssd2 vssd2 vccd2 vccd2 _7798_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_431 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_107_149 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_80_518 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6749_ _6749_/A _6749_/B vssd2 vssd2 vccd2 vccd2 _6750_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_456 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_478 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_103_366 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_103_399 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1541 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_515 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_113_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1585 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_161 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4713__A _4896_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_56_537 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_92 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_70 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_81 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5528__B _5528_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_98_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_64_592 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_3_306 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__3993__A_N _4267_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_51_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_456 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_51_286 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5080_ _5210_/B _5406_/A _5468_/A _5210_/A vssd2 vssd2 vccd2 vccd2 _5082_/A sky130_fd_sc_hd__o22ai_2
XFILLER_0_47_44 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4100_ _4656_/A _4100_/B vssd2 vssd2 vccd2 vccd2 _4101_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_66 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__3999__A _7763_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4031_ _4814_/B _4252_/D _4063_/B vssd2 vssd2 vccd2 vccd2 _4032_/C sky130_fd_sc_hd__and3_1
XFILLER_0_47_99 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_78_117 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_63_10 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_78_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_63_54 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6785__A1 _7094_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5982_ _5975_/X _5977_/X _5980_/X _5981_/X _5811_/C vssd2 vssd2 vccd2 vccd2 _6738_/A
+ sky130_fd_sc_hd__o41a_4
X_4933_ _5011_/A _5076_/D vssd2 vssd2 vccd2 vccd2 _4935_/A sky130_fd_sc_hd__or2_1
XANTENNA__6785__B2 _7047_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7721_ _7758_/CLK _7721_/D vssd2 vssd2 vccd2 vccd2 _7721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4864_ _4864_/A _4864_/B vssd2 vssd2 vccd2 vccd2 _4874_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_74_345 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7652_ _7800_/CLK _7652_/D vssd2 vssd2 vccd2 vccd2 _7652_/Q sky130_fd_sc_hd__dfxtp_1
X_7583_ _7590_/A vssd2 vssd2 vccd2 vccd2 _7583_/Y sky130_fd_sc_hd__inv_2
X_6603_ _6603_/A _6603_/B vssd2 vssd2 vccd2 vccd2 _6604_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_4795_ _4805_/A vssd2 vssd2 vccd2 vccd2 _4795_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4342__B _4896_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3815_ _3822_/A _3822_/B _3822_/C _3888_/B vssd2 vssd2 vccd2 vccd2 _3819_/B sky130_fd_sc_hd__o31a_2
X_6534_ _6337_/A _6337_/B _6453_/B _6452_/B _6452_/A vssd2 vssd2 vccd2 vccd2 _6536_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_103_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_27_294 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6465_ _6466_/A _6465_/B vssd2 vssd2 vccd2 vccd2 _7819_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_478 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_113_653 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_112_141 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_70_595 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5454__A _5454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_30_415 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5416_ _5417_/A _5417_/B vssd2 vssd2 vccd2 vccd2 _5461_/B sky130_fd_sc_hd__or2_1
Xoutput120 hold641/X vssd2 vssd2 vccd2 vccd2 hold290/A sky130_fd_sc_hd__buf_6
Xoutput131 hold639/X vssd2 vssd2 vccd2 vccd2 hold288/A sky130_fd_sc_hd__buf_6
X_6396_ _6670_/A _6396_/B vssd2 vssd2 vccd2 vccd2 _6396_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
Xoutput142 _7712_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[17] sky130_fd_sc_hd__buf_12
X_5347_ _5347_/A _5347_/B vssd2 vssd2 vccd2 vccd2 _5349_/B sky130_fd_sc_hd__xor2_1
Xoutput153 _7722_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[27] sky130_fd_sc_hd__buf_12
Xoutput164 _7703_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[8] sky130_fd_sc_hd__buf_12
X_5278_ _5279_/A _5279_/B vssd2 vssd2 vccd2 vccd2 _5313_/A sky130_fd_sc_hd__nor2_1
X_7017_ _7017_/A _7017_/B vssd2 vssd2 vccd2 vccd2 _7019_/B sky130_fd_sc_hd__xnor2_1
X_4229_ _4229_/A _4229_/B _4230_/B vssd2 vssd2 vccd2 vccd2 _4260_/A sky130_fd_sc_hd__and3_1
XFILLER_0_69_117 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6225__B1 _6152_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_437 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_84_109 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_93_643 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_93_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_92_153 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_53_529 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_18_261 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_92_197 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5364__A _5414_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5083__B _5431_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_108_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4708__A _4708_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_17_36 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7008__A2 _7255_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6923__A _7037_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_75_109 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_69_673 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_96_481 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__6642__B _6642_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_68_161 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_29_526 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_33_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_33_68 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1393 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_654 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_83_131 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_68_194 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_71_315 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_71_304 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7176__D _7253_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_37_570 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_114_417 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4580_ _4580_/A _4580_/B vssd2 vssd2 vccd2 vccd2 _4581_/B sky130_fd_sc_hd__xnor2_2
Xinput11 input11/A vssd2 vssd2 vccd2 vccd2 input11/X sky130_fd_sc_hd__clkbuf_1
Xinput22 input22/A vssd2 vssd2 vccd2 vccd2 input22/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xinput33 input33/A vssd2 vssd2 vccd2 vccd2 input33/X sky130_fd_sc_hd__clkbuf_1
Xinput44 input44/A vssd2 vssd2 vccd2 vccd2 input44/X sky130_fd_sc_hd__clkbuf_1
Xinput55 wbs_adr_i[14] vssd2 vssd2 vccd2 vccd2 _7343_/D sky130_fd_sc_hd__clkbuf_1
Xinput88 input88/A vssd2 vssd2 vccd2 vccd2 input88/X sky130_fd_sc_hd__clkbuf_1
Xinput66 wbs_adr_i[24] vssd2 vssd2 vccd2 vccd2 _7339_/B sky130_fd_sc_hd__clkbuf_1
Xinput77 wbs_adr_i[5] vssd2 vssd2 vccd2 vccd2 _7342_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__6089__B _6783_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6250_ _6250_/A _6316_/B vssd2 vssd2 vccd2 vccd2 _7816_/D sky130_fd_sc_hd__xnor2_1
Xinput99 wbs_stb_i vssd2 vssd2 vccd2 vccd2 _7453_/B sky130_fd_sc_hd__clkbuf_2
X_6181_ _6182_/A _6182_/B vssd2 vssd2 vccd2 vccd2 _6181_/Y sky130_fd_sc_hd__nand2_1
X_5201_ _5201_/A _5201_/B _5201_/C vssd2 vssd2 vccd2 vccd2 _5201_/X sky130_fd_sc_hd__and3_1
X_5132_ _5133_/D _5132_/B vssd2 vssd2 vccd2 vccd2 _7745_/D sky130_fd_sc_hd__xor2_1
XANTENNA__5721__B _5781_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5063_ _5063_/A _5063_/B vssd2 vssd2 vccd2 vccd2 _5064_/B sky130_fd_sc_hd__xor2_4
X_4014_ _4002_/Y _4004_/Y _4086_/B _3893_/B _3994_/X vssd2 vssd2 vccd2 vccd2 _4014_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_90_41 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_87_492 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5965_ _5965_/A _5969_/A vssd2 vssd2 vccd2 vccd2 _5966_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_610 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_47_323 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_90_85 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4916_ _4916_/A _4916_/B vssd2 vssd2 vccd2 vccd2 _4919_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_131 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7704_ _7802_/CLK _7704_/D vssd2 vssd2 vccd2 vccd2 _7704_/Q sky130_fd_sc_hd__dfxtp_1
X_5896_ _5713_/Y _5896_/B vssd2 vssd2 vccd2 vccd2 _5896_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_0_114_81 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_90_602 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_74_153 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_62_304 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__5168__B _5528_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4847_ _5455_/A _4847_/B vssd2 vssd2 vccd2 vccd2 _4848_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_442 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7635_ _7641_/A vssd2 vssd2 vccd2 vccd2 _7635_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_105_417 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_74_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_7_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_15_220 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_90_668 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4778_ _4778_/A _4778_/B vssd2 vssd2 vccd2 vccd2 _4780_/A sky130_fd_sc_hd__nand2_2
X_7566_ _7613_/A vssd2 vssd2 vccd2 vccd2 _7566_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_540 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_7_486 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6517_ _6668_/A _6430_/B _6438_/B _6436_/X vssd2 vssd2 vccd2 vccd2 _6519_/B sky130_fd_sc_hd__a31o_1
XANTENNA__4800__B _5030_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7497_ _7524_/A vssd2 vssd2 vccd2 vccd2 _7497_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_264 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_30_212 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_113_461 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6448_ _6449_/A _6449_/B vssd2 vssd2 vccd2 vccd2 _6448_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_70_392 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7486__A2 _7453_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6379_ _6380_/A _6380_/B vssd2 vssd2 vccd2 vccd2 _6379_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_100_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5497__B2 _5498_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5497__A1 _5550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_30_267 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_100_177 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4528__A _4962_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5359__A _5454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_93_440 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5972__A2 _5786_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_108_233 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_93_484 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_81_602 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5078__B _5145_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_65_164 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_65_142 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7574__A _7613_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_53_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_108_277 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_80_145 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_34_573 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_4_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7854_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__7477__A2 _7483_/A2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_418 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_46 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_44_23 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_88_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_44_45 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_88_289 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_76_429 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_44_89 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5750_ _7840_/Q _6510_/B vssd2 vssd2 vccd2 vccd2 _5750_/X sky130_fd_sc_hd__and2_1
XFILLER_0_29_323 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_29_345 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4173__A _4598_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4701_ _4699_/A _4631_/B _4640_/B _4638_/X vssd2 vssd2 vccd2 vccd2 _4722_/A sky130_fd_sc_hd__a31oi_2
XTAP_1190 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5681_ _7880_/Q _5681_/B vssd2 vssd2 vccd2 vccd2 _6152_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_84_484 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4632_ _4704_/B _5276_/A vssd2 vssd2 vccd2 vccd2 _4636_/A sky130_fd_sc_hd__or2_1
XFILLER_0_56_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_44_326 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7420_ _7420_/A _7420_/B vssd2 vssd2 vccd2 vccd2 _7451_/S sky130_fd_sc_hd__or2_4
XFILLER_0_114_225 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_71_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_4_412 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4563_ _4966_/A _4711_/A _4782_/B _4896_/A vssd2 vssd2 vccd2 vccd2 _4565_/A sky130_fd_sc_hd__o22ai_1
XFILLER_0_69_20 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7351_ _7387_/A _7386_/A hold99/X vssd2 vssd2 vccd2 vccd2 _7351_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_4_467 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold603 hold96/X vssd2 vssd2 vccd2 vccd2 _7871_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 hold625/A vssd2 vssd2 vccd2 vccd2 hold625/X sky130_fd_sc_hd__dlygate4sd3_1
X_6302_ _6302_/A _6302_/B vssd2 vssd2 vccd2 vccd2 _6303_/B sky130_fd_sc_hd__xnor2_2
Xhold636 _7825_/Q vssd2 vssd2 vccd2 vccd2 hold636/X sky130_fd_sc_hd__dlygate4sd3_1
X_7282_ _7283_/B _7283_/C _7283_/A vssd2 vssd2 vccd2 vccd2 _7308_/B sky130_fd_sc_hd__a21o_2
X_4494_ _4898_/A _5276_/A vssd2 vssd2 vccd2 vccd2 _4498_/A sky130_fd_sc_hd__nor2_1
Xhold614 _7808_/Q vssd2 vssd2 vccd2 vccd2 hold614/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7468__A2 _7483_/A2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold669 hold669/A vssd2 vssd2 vccd2 vccd2 hold669/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 _7830_/Q vssd2 vssd2 vccd2 vccd2 hold658/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold647 hold647/A vssd2 vssd2 vccd2 vccd2 hold647/X sky130_fd_sc_hd__dlygate4sd3_1
X_6233_ _6233_/A _6233_/B vssd2 vssd2 vccd2 vccd2 _6234_/B sky130_fd_sc_hd__xor2_1
XANTENNA__7423__S _7451_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6164_ _6164_/A _6164_/B vssd2 vssd2 vccd2 vccd2 _6165_/B sky130_fd_sc_hd__xnor2_2
XTAP_952 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _5115_/A _5115_/B vssd2 vssd2 vccd2 vccd2 _5118_/A sky130_fd_sc_hd__xnor2_4
XTAP_996 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _5691_/A _5691_/B _6094_/B _6155_/B _6358_/A vssd2 vssd2 vccd2 vccd2 _6095_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__5451__B _5451_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_fanout191_A _5366_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_109_81 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5046_ _5047_/A _5047_/B vssd2 vssd2 vccd2 vccd2 _5046_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout289_A _7629_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_33_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__4067__B _4893_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5403__A1 _5498_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6997_ _6997_/A _6997_/B vssd2 vssd2 vccd2 vccd2 _6999_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__7097__C _7222_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5948_ _5945_/X _5947_/X _5755_/C vssd2 vssd2 vccd2 vccd2 _5948_/X sky130_fd_sc_hd__o21a_4
XANTENNA__5403__B2 _5404_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4083__A _7763_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5954__A2 _6150_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_48_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_90_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5879_ _6282_/A _6071_/B _6019_/C _6019_/D vssd2 vssd2 vccd2 vccd2 _5886_/B sky130_fd_sc_hd__and4_1
XFILLER_0_35_326 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_105_225 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_50_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7618_ _7645_/A vssd2 vssd2 vccd2 vccd2 _7618_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5167__B1 _5374_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7549_ _7565_/A vssd2 vssd2 vccd2 vccd2 _7549_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7459__A2 _7454_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6738__A _6738_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5642__A _6424_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_101_497 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_101_486 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4258__A _4598_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7569__A _7613_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_105_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_98_587 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_14_48 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_26_304 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_93_281 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_38_175 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_38_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_26_348 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_81_498 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_81_487 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_111_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4381__A1 _7772_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4381__B2 _4809_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_237 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4168__A _7765_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3800__A _6253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6920_ _6073_/Y _6920_/A2 _7291_/A _5664_/C vssd2 vssd2 vccd2 vccd2 _6922_/A sky130_fd_sc_hd__a211o_1
XFILLER_0_76_204 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_71_10 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6851_ _5991_/X _5993_/X _7222_/C _5781_/B vssd2 vssd2 vccd2 vccd2 _6854_/A sky130_fd_sc_hd__o211a_1
XFILLER_0_49_418 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_76_259 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_71_54 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5802_ _6398_/A _5836_/B _5665_/B _6283_/A _5878_/B vssd2 vssd2 vccd2 vccd2 _5803_/D
+ sky130_fd_sc_hd__a32o_1
X_6782_ _6782_/A _6782_/B vssd2 vssd2 vccd2 vccd2 _6784_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_473 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_9_537 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3994_ _4457_/A _4458_/C _4141_/C _4082_/D vssd2 vssd2 vccd2 vccd2 _3994_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_44_123 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5733_ _7873_/Q _5734_/B vssd2 vssd2 vccd2 vccd2 _5762_/B sky130_fd_sc_hd__xor2_1
XANTENNA__7418__S _7418_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5664_ _6157_/A _7855_/Q _5664_/C _5811_/B vssd2 vssd2 vccd2 vccd2 _5664_/X sky130_fd_sc_hd__and4_1
X_4615_ _4543_/A _4543_/B _4541_/X vssd2 vssd2 vccd2 vccd2 _4617_/B sky130_fd_sc_hd__a21oi_2
X_7403_ _7440_/A _7403_/B vssd2 vssd2 vccd2 vccd2 _7670_/D sky130_fd_sc_hd__and2_1
XFILLER_0_25_370 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_32_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5595_ _7868_/Q _5598_/B vssd2 vssd2 vccd2 vccd2 _5659_/A sky130_fd_sc_hd__xor2_1
X_7334_ _7334_/A _7334_/B _7334_/C _7334_/D vssd2 vssd2 vccd2 vccd2 _7334_/X sky130_fd_sc_hd__and4_1
Xhold400 hold696/X vssd2 vssd2 vccd2 vccd2 _7801_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 _7775_/Q vssd2 vssd2 vccd2 vccd2 hold411/X sky130_fd_sc_hd__dlygate4sd3_1
X_4546_ _4547_/A _4547_/B vssd2 vssd2 vccd2 vccd2 _4619_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_111_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold422 input36/X vssd2 vssd2 vccd2 vccd2 hold2/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 hold33/X vssd2 vssd2 vccd2 vccd2 input31/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 la_data_in[12] vssd2 vssd2 vccd2 vccd2 hold17/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_351 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold455 hold26/X vssd2 vssd2 vccd2 vccd2 _7853_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7265_ _7263_/Y _7264_/Y _7224_/A _7291_/B vssd2 vssd2 vccd2 vccd2 _7267_/B sky130_fd_sc_hd__o2bb2a_1
Xhold466 input35/X vssd2 vssd2 vccd2 vccd2 hold24/A sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap185 _5984_/B vssd2 vssd2 vccd2 vccd2 _6873_/A sky130_fd_sc_hd__clkbuf_2
Xhold477 hold13/X vssd2 vssd2 vccd2 vccd2 input13/A sky130_fd_sc_hd__dlygate4sd3_1
X_4477_ _4478_/A _4478_/B vssd2 vssd2 vccd2 vccd2 _4547_/A sky130_fd_sc_hd__nor2_1
X_6216_ _6216_/A _6216_/B vssd2 vssd2 vccd2 vccd2 _6217_/B sky130_fd_sc_hd__nand2_1
X_7196_ _7196_/A _7196_/B vssd2 vssd2 vccd2 vccd2 _7199_/B sky130_fd_sc_hd__xnor2_1
Xhold499 hold52/X vssd2 vssd2 vccd2 vccd2 _7856_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 la_data_in[15] vssd2 vssd2 vccd2 vccd2 hold27/A sky130_fd_sc_hd__dlygate4sd3_1
X_6147_ _6812_/A _6812_/B _6705_/B _6939_/A vssd2 vssd2 vccd2 vccd2 _6148_/B sky130_fd_sc_hd__or4_1
XTAP_760 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__7389__A _7440_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6078_ _6078_/A _6078_/B _6078_/C _6078_/D vssd2 vssd2 vccd2 vccd2 _6078_/Y sky130_fd_sc_hd__nor4_1
X_5029_ _5029_/A _5498_/D vssd2 vssd2 vccd2 vccd2 _5029_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_218 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_48_440 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_75_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_90_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_106_567 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_63_487 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_31_362 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6104__A2 _6150_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_101_261 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_98_362 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_86_524 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_86_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6634__C _7222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_73_218 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__6040__A1 _6283_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_73_229 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_26_101 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_109_361 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_54_454 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_26_145 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_81_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4400_ _4882_/A _5099_/A _4401_/A vssd2 vssd2 vccd2 vccd2 _4400_/X sky130_fd_sc_hd__or3_1
XFILLER_0_41_126 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5380_ _5412_/A _5380_/B vssd2 vssd2 vccd2 vccd2 _5381_/B sky130_fd_sc_hd__nor2_1
X_4331_ _4809_/A _4082_/B _4328_/X _4330_/X vssd2 vssd2 vccd2 vccd2 _4331_/X sky130_fd_sc_hd__a211o_2
XFILLER_0_10_524 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_22_373 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7050_ _7143_/A _7222_/B vssd2 vssd2 vccd2 vccd2 _7052_/B sky130_fd_sc_hd__nand2_1
Xfanout209 _4807_/A vssd2 vssd2 vccd2 vccd2 _4962_/A sky130_fd_sc_hd__buf_4
X_4262_ _7768_/Q _4454_/B vssd2 vssd2 vccd2 vccd2 _4262_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4106__A1 _7763_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4106__B2 _7764_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6001_ _6001_/A _6001_/B _6001_/C vssd2 vssd2 vccd2 vccd2 _6003_/B sky130_fd_sc_hd__nand3_2
XANTENNA__4657__A2 _5458_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4193_ _4193_/A _4193_/B vssd2 vssd2 vccd2 vccd2 _4196_/B sky130_fd_sc_hd__nor2_1
X_6903_ _6904_/B _6904_/A vssd2 vssd2 vccd2 vccd2 _6903_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_77_513 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_49_237 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7883_ _7886_/CLK _7883_/D _7642_/Y vssd2 vssd2 vccd2 vccd2 _7883_/Q sky130_fd_sc_hd__dfrtp_4
X_6834_ _6834_/A _6834_/B vssd2 vssd2 vccd2 vccd2 _6839_/B sky130_fd_sc_hd__xor2_2
X_6765_ _6765_/A _6765_/B _6765_/C vssd2 vssd2 vccd2 vccd2 _6767_/B sky130_fd_sc_hd__or3_2
XFILLER_0_92_527 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3977_ _7760_/Q _4068_/B vssd2 vssd2 vccd2 vccd2 _3977_/X sky130_fd_sc_hd__and2_1
X_5716_ _7847_/Q _6155_/B _5769_/B _5944_/C vssd2 vssd2 vccd2 vccd2 _5716_/X sky130_fd_sc_hd__and4_1
X_6696_ _6696_/A _6769_/C vssd2 vssd2 vccd2 vccd2 _7822_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_498 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_32_104 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_60_446 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5647_ _7856_/Q _5647_/B vssd2 vssd2 vccd2 vccd2 _5812_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_137 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_103_548 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5578_ _7861_/Q _7862_/Q vssd2 vssd2 vccd2 vccd2 _5581_/C sky130_fd_sc_hd__or2_2
X_4529_ _4527_/X _4529_/B vssd2 vssd2 vccd2 vccd2 _4530_/B sky130_fd_sc_hd__and2b_1
X_7317_ _7263_/Y _7302_/B _7301_/A vssd2 vssd2 vccd2 vccd2 _7319_/C sky130_fd_sc_hd__o21a_1
Xhold252 _7456_/X vssd2 vssd2 vccd2 vccd2 _7696_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 _7731_/Q vssd2 vssd2 vccd2 vccd2 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 _7465_/X vssd2 vssd2 vccd2 vccd2 _7705_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_170 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
Xhold285 hold642/X vssd2 vssd2 vccd2 vccd2 hold643/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 hold274/A vssd2 vssd2 vccd2 vccd2 la_data_out[21] sky130_fd_sc_hd__buf_12
X_7248_ _7279_/A _7217_/B _7210_/A vssd2 vssd2 vccd2 vccd2 _7249_/B sky130_fd_sc_hd__a21bo_1
Xhold296 hold296/A vssd2 vssd2 vccd2 vccd2 la_data_out[12] sky130_fd_sc_hd__buf_12
Xhold263 hold616/X vssd2 vssd2 vccd2 vccd2 hold617/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_192 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7179_ _7179_/A _7179_/B vssd2 vssd2 vccd2 vccd2 _7188_/A sky130_fd_sc_hd__xnor2_1
XTAP_590 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5073__A2 _5431_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_95_376 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_83_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_36_421 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_102_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_51_402 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_36_465 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_23_137 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_36_498 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_23_159 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_592 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_36_35 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_36_46 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
Xinput9 input9/A vssd2 vssd2 vccd2 vccd2 input9/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3988__C _4656_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_36_68 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_86_376 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6013__A1 _6402_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4880_ _5029_/A _4880_/B vssd2 vssd2 vccd2 vccd2 _4883_/A sky130_fd_sc_hd__or2_1
X_3900_ _3886_/X _3899_/X _3898_/X _3892_/X vssd2 vssd2 vccd2 vccd2 _3900_/X sky130_fd_sc_hd__a211o_1
X_3831_ _7801_/Q _3831_/B vssd2 vssd2 vccd2 vccd2 _3886_/C sky130_fd_sc_hd__xnor2_2
X_6550_ _6550_/A _7255_/B vssd2 vssd2 vccd2 vccd2 _6551_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_39_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5501_ _5470_/A _5470_/B _5466_/A vssd2 vssd2 vccd2 vccd2 _5503_/B sky130_fd_sc_hd__o21a_1
X_6481_ _6481_/A _6481_/B _6481_/C vssd2 vssd2 vccd2 vccd2 _6483_/A sky130_fd_sc_hd__and3_1
XFILLER_0_112_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4327__A1 _7772_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5432_ _5433_/B _5433_/C _5433_/A vssd2 vssd2 vccd2 vccd2 _5480_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_112_345 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_23_671 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5363_ _5363_/A _5363_/B vssd2 vssd2 vccd2 vccd2 _5365_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_112_389 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7102_ _7103_/A _7103_/B vssd2 vssd2 vccd2 vccd2 _7102_/Y sky130_fd_sc_hd__nand2b_1
X_4314_ _4125_/C _4311_/X _4313_/X vssd2 vssd2 vccd2 vccd2 _4314_/X sky130_fd_sc_hd__a21o_1
X_5294_ _5295_/A _5295_/B _5293_/Y vssd2 vssd2 vccd2 vccd2 _5294_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_10_376 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5827__A1 _6282_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7033_ _7033_/A _7033_/B _7033_/C _7033_/D vssd2 vssd2 vccd2 vccd2 _7326_/A sky130_fd_sc_hd__and4_2
X_4245_ _4303_/B _4303_/C vssd2 vssd2 vccd2 vccd2 _4247_/B sky130_fd_sc_hd__or2_1
XANTENNA__7431__S _7451_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4176_ _4177_/A _4177_/B vssd2 vssd2 vccd2 vccd2 _4176_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6252__A1 _7850_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6252__B2 _6283_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_89_181 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1019 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_365 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6571__A _6571_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7866_ _7870_/CLK _7866_/D _7625_/Y vssd2 vssd2 vccd2 vccd2 _7866_/Q sky130_fd_sc_hd__dfrtp_4
X_6817_ _6742_/A _6741_/B _6741_/A vssd2 vssd2 vccd2 vccd2 _6819_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_9_131 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7797_ _7798_/CLK _7797_/D _7556_/Y vssd2 vssd2 vccd2 vccd2 _7797_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_443 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6748_ _6749_/A _6749_/B vssd2 vssd2 vccd2 vccd2 _6748_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_45_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_413 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6679_ _6680_/A _6680_/B vssd2 vssd2 vccd2 vccd2 _6679_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_5_370 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_378 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_13_192 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_96_641 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1542 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_549 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XPHY_60 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_71 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_82 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4713__B _5276_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XPHY_93 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_64_571 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_36_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_20_641 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5809__A1 _7850_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4030_ _4252_/B _4030_/B _4427_/A vssd2 vssd2 vccd2 vccd2 _4030_/X sky130_fd_sc_hd__and3_2
XFILLER_0_99_490 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6785__A2 _7143_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5981_ _6157_/A _5810_/X _6017_/B _7847_/Q _5978_/X vssd2 vssd2 vccd2 vccd2 _5981_/X
+ sky130_fd_sc_hd__a221o_1
X_4932_ _4874_/A _4874_/B _4873_/A vssd2 vssd2 vccd2 vccd2 _4951_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_47_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7720_ _7723_/CLK _7720_/D vssd2 vssd2 vccd2 vccd2 _7720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_313 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_47_516 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7651_ _7779_/CLK _7651_/D vssd2 vssd2 vccd2 vccd2 _7651_/Q sky130_fd_sc_hd__dfxtp_1
X_6602_ _6603_/A _6603_/B vssd2 vssd2 vccd2 vccd2 _6602_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_86_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4863_ _4863_/A _5550_/A vssd2 vssd2 vccd2 vccd2 _4864_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_74_357 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_6_101 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7582_ _7590_/A vssd2 vssd2 vccd2 vccd2 _7582_/Y sky130_fd_sc_hd__inv_2
X_4794_ _4730_/A _4730_/B _4727_/Y vssd2 vssd2 vccd2 vccd2 _4805_/A sky130_fd_sc_hd__o21ai_4
X_3814_ _7799_/Q _7800_/Q _7801_/Q _7802_/Q vssd2 vssd2 vccd2 vccd2 _3822_/C sky130_fd_sc_hd__or4_2
XANTENNA__6942__C1 _7143_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6533_ _6533_/A _6533_/B vssd2 vssd2 vccd2 vccd2 _6536_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_109 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_82_390 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6464_ _7336_/A _6466_/B vssd2 vssd2 vccd2 vccd2 _6465_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_70_552 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_113_665 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xoutput110 hold637/X vssd2 vssd2 vccd2 vccd2 hold284/A sky130_fd_sc_hd__buf_6
XFILLER_0_88_41 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5415_ _5415_/A _5462_/A vssd2 vssd2 vccd2 vccd2 _5417_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_113_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xoutput121 hold669/X vssd2 vssd2 vccd2 vccd2 hold316/A sky130_fd_sc_hd__buf_6
XFILLER_0_112_153 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6395_ _6348_/A _6348_/B _6346_/X vssd2 vssd2 vccd2 vccd2 _6411_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_88_85 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xoutput132 hold631/X vssd2 vssd2 vccd2 vccd2 hold280/A sky130_fd_sc_hd__buf_6
Xoutput143 _7713_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[18] sky130_fd_sc_hd__buf_12
XFILLER_0_112_197 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5346_ _5347_/B _5347_/A vssd2 vssd2 vccd2 vccd2 _5395_/A sky130_fd_sc_hd__nand2b_1
Xoutput165 _7704_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[9] sky130_fd_sc_hd__buf_12
Xoutput154 _7723_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[28] sky130_fd_sc_hd__buf_12
X_5277_ _5210_/B _5498_/D _5550_/B _5210_/A vssd2 vssd2 vccd2 vccd2 _5279_/B sky130_fd_sc_hd__o22a_1
X_7016_ _7017_/A _7017_/B vssd2 vssd2 vccd2 vccd2 _7081_/A sky130_fd_sc_hd__nor2_1
X_4228_ _4228_/A _4228_/B vssd2 vssd2 vccd2 vccd2 _4230_/B sky130_fd_sc_hd__xnor2_1
X_4159_ _4454_/A _4251_/B vssd2 vssd2 vccd2 vccd2 _4171_/A sky130_fd_sc_hd__and2_1
XFILLER_0_97_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__7397__A _7440_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_38_516 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_92_121 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7849_ _7854_/CLK _7849_/D _7608_/Y vssd2 vssd2 vccd2 vccd2 _7849_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_92_165 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_18_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_243 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_104_654 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_585 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_21_405 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5364__B _5550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_104_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_21_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4708__B _5550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6923__B _7224_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_641 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_96_471 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1350 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_96_493 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1383 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__3985__D _5030_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1394 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 input12/A vssd2 vssd2 vccd2 vccd2 input12/X sky130_fd_sc_hd__clkbuf_1
Xinput45 input45/A vssd2 vssd2 vccd2 vccd2 input45/X sky130_fd_sc_hd__clkbuf_1
Xinput23 input23/A vssd2 vssd2 vccd2 vccd2 input23/X sky130_fd_sc_hd__clkbuf_1
Xinput34 input34/A vssd2 vssd2 vccd2 vccd2 input34/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_416 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xinput56 wbs_adr_i[15] vssd2 vssd2 vccd2 vccd2 _7343_/C sky130_fd_sc_hd__clkbuf_1
Xinput89 input89/A vssd2 vssd2 vccd2 vccd2 input89/X sky130_fd_sc_hd__clkbuf_1
Xinput78 wbs_adr_i[6] vssd2 vssd2 vccd2 vccd2 _7342_/D sky130_fd_sc_hd__buf_1
Xinput67 wbs_adr_i[25] vssd2 vssd2 vccd2 vccd2 _7339_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_159 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6089__C _6812_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6180_ _6180_/A _6180_/B vssd2 vssd2 vccd2 vccd2 _6182_/B sky130_fd_sc_hd__xnor2_2
X_5200_ _5201_/A _5201_/B _5201_/C vssd2 vssd2 vccd2 vccd2 _5301_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_20_460 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_58_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5131_ _5133_/A _5133_/B _5133_/C _5548_/A vssd2 vssd2 vccd2 vccd2 _5132_/B sky130_fd_sc_hd__a31o_1
X_5062_ _5063_/A _5063_/B vssd2 vssd2 vccd2 vccd2 _5062_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3803__A _7842_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4013_ _3999_/Y _4011_/Y _4012_/Y _3893_/D vssd2 vssd2 vccd2 vccd2 _4017_/A sky130_fd_sc_hd__a31o_1
XANTENNA__4634__A _4966_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_94_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_90_53 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5964_ _5965_/A _5969_/A vssd2 vssd2 vccd2 vccd2 _6064_/A sky130_fd_sc_hd__or2_1
XFILLER_0_47_313 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7703_ _7798_/CLK _7703_/D vssd2 vssd2 vccd2 vccd2 _7703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_97 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4915_ _4915_/A _4915_/B vssd2 vssd2 vccd2 vccd2 _4916_/B sky130_fd_sc_hd__xor2_4
X_5895_ _5755_/C _5853_/B _5894_/X _6094_/B _7845_/Q vssd2 vssd2 vccd2 vccd2 _5896_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_74_165 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4846_ _4769_/B _4849_/C vssd2 vssd2 vccd2 vccd2 _4847_/B sky130_fd_sc_hd__nand2b_1
X_7634_ _7641_/A vssd2 vssd2 vccd2 vccd2 _7634_/Y sky130_fd_sc_hd__inv_2
X_7565_ _7565_/A vssd2 vssd2 vccd2 vccd2 _7565_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_465 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_105_429 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_99_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4777_ _4863_/A _5011_/A _5142_/C _5076_/D vssd2 vssd2 vccd2 vccd2 _4778_/B sky130_fd_sc_hd__or4_1
X_6516_ _6516_/A _6516_/B vssd2 vssd2 vccd2 vccd2 _6519_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__4800__C _4800_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7496_ _7524_/A vssd2 vssd2 vccd2 vccd2 _7496_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_113_473 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6447_ _6373_/A _6373_/B _6371_/Y vssd2 vssd2 vccd2 vccd2 _6449_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_30_224 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6378_ _6303_/A _6303_/B _6301_/X vssd2 vssd2 vccd2 vccd2 _6380_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__5497__A2 _5528_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_30_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5329_ _5329_/A _5329_/B vssd2 vssd2 vccd2 vccd2 _5330_/B sky130_fd_sc_hd__and2_1
XFILLER_0_100_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4809__A _4809_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4528__B _4966_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_78_482 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_93_430 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_38_346 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_108_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_93_496 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_108_289 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_419 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7740__D _7740_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_57_600 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4454__A _4454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_493 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XTAP_1191 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _4839_/A _4700_/B vssd2 vssd2 vccd2 vccd2 _4762_/A sky130_fd_sc_hd__and2_1
XFILLER_0_56_165 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5680_ _7879_/Q _5694_/A _5694_/B _5694_/C _5735_/B vssd2 vssd2 vccd2 vccd2 _5681_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_0_29_379 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4631_ _4699_/A _4631_/B vssd2 vssd2 vccd2 vccd2 _4640_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5285__A _5328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_37_390 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_114_237 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4562_ _4736_/A _5276_/A vssd2 vssd2 vccd2 vccd2 _4566_/A sky130_fd_sc_hd__or2_1
XFILLER_0_71_179 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7350_ _7453_/C _7453_/B _7350_/C vssd2 vssd2 vccd2 vccd2 _7387_/A sky130_fd_sc_hd__nand3_1
X_6301_ _6302_/A _6302_/B vssd2 vssd2 vccd2 vccd2 _6301_/X sky130_fd_sc_hd__and2b_1
Xhold626 _7826_/Q vssd2 vssd2 vccd2 vccd2 hold626/X sky130_fd_sc_hd__dlygate4sd3_1
X_7281_ _7210_/A _7247_/A _7247_/B vssd2 vssd2 vccd2 vccd2 _7283_/C sky130_fd_sc_hd__a21bo_1
Xhold615 hold615/A vssd2 vssd2 vccd2 vccd2 hold615/X sky130_fd_sc_hd__dlygate4sd3_1
X_4493_ _4598_/A _5142_/C vssd2 vssd2 vccd2 vccd2 _4502_/A sky130_fd_sc_hd__or2_1
Xhold604 la_data_in[2] vssd2 vssd2 vccd2 vccd2 hold93/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_110_421 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold659 hold659/A vssd2 vssd2 vccd2 vccd2 hold659/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold637 hold637/A vssd2 vssd2 vccd2 vccd2 hold637/X sky130_fd_sc_hd__dlygate4sd3_1
X_6232_ _6233_/A _6233_/B vssd2 vssd2 vccd2 vccd2 _6232_/Y sky130_fd_sc_hd__nor2_1
Xhold648 _7819_/Q vssd2 vssd2 vccd2 vccd2 hold648/X sky130_fd_sc_hd__dlygate4sd3_1
X_6163_ _6590_/A _6164_/A _7094_/A vssd2 vssd2 vccd2 vccd2 _6163_/X sky130_fd_sc_hd__and3_1
XANTENNA__6428__A1 _6738_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4629__A _4708_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_953 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5114_/A _5114_/B vssd2 vssd2 vccd2 vccd2 _5115_/B sky130_fd_sc_hd__xnor2_4
XTAP_986 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6158_/A _6094_/B vssd2 vssd2 vccd2 vccd2 _6094_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_109_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_997 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5220_/A _4965_/B _4970_/B _4968_/Y vssd2 vssd2 vccd2 vccd2 _5047_/B sky130_fd_sc_hd__o31a_2
XFILLER_0_79_202 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_26_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_79_235 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_79_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6996_ _7140_/A _7181_/A vssd2 vssd2 vccd2 vccd2 _6997_/B sky130_fd_sc_hd__nor2_1
XANTENNA__7097__D _7294_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5947_ _5947_/A _5947_/B _5947_/C _5947_/D vssd2 vssd2 vccd2 vccd2 _5947_/X sky130_fd_sc_hd__or4_4
XANTENNA__5403__A2 _5468_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_90_433 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_75_496 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5907__B _6634_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_62_102 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5878_ _6398_/A _5878_/B _5878_/C vssd2 vssd2 vccd2 vccd2 _5883_/C sky130_fd_sc_hd__and3_1
XANTENNA__5757__A_N _5992_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7617_ _7645_/A vssd2 vssd2 vccd2 vccd2 _7617_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_90_455 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4829_ _4829_/A _4829_/B vssd2 vssd2 vccd2 vccd2 _4830_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_62_157 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_105_237 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_90_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7548_ _7564_/A vssd2 vssd2 vccd2 vccd2 _7548_/Y sky130_fd_sc_hd__inv_2
X_7479_ _7719_/Q _7483_/A2 _7483_/B1 hold339/X vssd2 vssd2 vccd2 vccd2 _7479_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_113_281 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6738__B _7099_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4258__B _4711_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_58_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_78_290 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_66_452 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_81_433 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_53_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_93_293 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_81_444 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_81_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_22_500 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_22_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA_max_cap247_A _4006_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_39_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_238 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6664__A _6664_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold1 hold1/A vssd2 vssd2 vccd2 vccd2 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_522 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5094__B1 _5550_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_89_588 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6850_ _6808_/A _6808_/C _6808_/B vssd2 vssd2 vccd2 vccd2 _6868_/A sky130_fd_sc_hd__a21boi_1
X_6781_ _6855_/A _6939_/A _7253_/A _7253_/B vssd2 vssd2 vccd2 vccd2 _6782_/B sky130_fd_sc_hd__or4_1
X_5801_ _5607_/A _5607_/B _5620_/B _5620_/C _5653_/C vssd2 vssd2 vccd2 vccd2 _6075_/D
+ sky130_fd_sc_hd__o2111a_2
X_5732_ _5739_/A _5755_/C vssd2 vssd2 vccd2 vccd2 _5853_/A sky130_fd_sc_hd__nor2_1
X_3993_ _4267_/D _3895_/C _4148_/B _3993_/D vssd2 vssd2 vccd2 vccd2 _4082_/D sky130_fd_sc_hd__and4bb_1
XFILLER_0_72_400 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_44_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_29_165 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5663_ _6071_/B _5921_/D vssd2 vssd2 vccd2 vccd2 _5663_/X sky130_fd_sc_hd__and2_1
XFILLER_0_72_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_60_617 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4614_ _4614_/A _4614_/B vssd2 vssd2 vccd2 vccd2 _4617_/A sky130_fd_sc_hd__xnor2_2
X_5594_ _7841_/Q _5594_/B _5594_/C vssd2 vssd2 vccd2 vccd2 _5594_/X sky130_fd_sc_hd__and3_1
X_7402_ hold139/X _7782_/D _7418_/S vssd2 vssd2 vccd2 vccd2 _7402_/X sky130_fd_sc_hd__mux2_1
X_7333_ _7333_/A _7333_/B vssd2 vssd2 vccd2 vccd2 _7836_/D sky130_fd_sc_hd__xnor2_1
X_4545_ _4545_/A _4545_/B vssd2 vssd2 vccd2 vccd2 _4547_/B sky130_fd_sc_hd__xnor2_2
Xhold401 _7661_/Q vssd2 vssd2 vccd2 vccd2 hold401/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold423 hold2/X vssd2 vssd2 vccd2 vccd2 _7848_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 input31/X vssd2 vssd2 vccd2 vccd2 hold34/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 hold17/X vssd2 vssd2 vccd2 vccd2 input4/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 _7805_/Q vssd2 vssd2 vccd2 vccd2 _3826_/A sky130_fd_sc_hd__buf_1
XFILLER_0_96_41 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7264_ _7264_/A _7264_/B vssd2 vssd2 vccd2 vccd2 _7264_/Y sky130_fd_sc_hd__nand2_1
Xhold467 hold24/X vssd2 vssd2 vccd2 vccd2 _7847_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 la_data_in[34] vssd2 vssd2 vccd2 vccd2 hold15/A sky130_fd_sc_hd__dlygate4sd3_1
X_4476_ _4413_/A _4413_/B _4411_/Y vssd2 vssd2 vccd2 vccd2 _4478_/B sky130_fd_sc_hd__a21boi_2
Xhold478 input13/X vssd2 vssd2 vccd2 vccd2 hold14/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_96_85 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6215_ _6812_/A _6812_/B _6215_/C _6989_/A vssd2 vssd2 vccd2 vccd2 _6216_/B sky130_fd_sc_hd__or4_1
X_7195_ _7196_/A _7196_/B vssd2 vssd2 vccd2 vccd2 _7244_/A sky130_fd_sc_hd__or2_1
Xhold489 hold27/X vssd2 vssd2 vccd2 vccd2 input7/A sky130_fd_sc_hd__dlygate4sd3_1
X_6146_ _6664_/A _5948_/X _5994_/X _5931_/C vssd2 vssd2 vccd2 vccd2 _6148_/A sky130_fd_sc_hd__a22o_1
XTAP_761 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _7847_/Q _7313_/A _6398_/B _7848_/Q vssd2 vssd2 vccd2 vccd2 _6078_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4806__B _5222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5028_ _5029_/A _5164_/B vssd2 vssd2 vccd2 vccd2 _5030_/D sky130_fd_sc_hd__nor2_1
X_6979_ _6979_/A _6979_/B vssd2 vssd2 vccd2 vccd2 _6979_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_422 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_48_474 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA_hold409_A _7806_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_8_582 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_579 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5653__A _7843_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_31_330 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_31_374 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_101_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6634__D _7222_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_58_205 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5828__A _7845_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_39_441 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_109_373 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_41_69 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_54_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_54_466 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_54_499 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5000__B1 _5548_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_41_149 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_105_590 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5551__A1 _4809_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4330_ _7771_/Q _3830_/X _4326_/D _4329_/X vssd2 vssd2 vccd2 vccd2 _4330_/X sky130_fd_sc_hd__a31o_1
X_4261_ _4356_/A _4261_/B vssd2 vssd2 vccd2 vccd2 _4294_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4106__A2 _4809_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6000_ _5952_/A _5952_/B _5952_/C vssd2 vssd2 vccd2 vccd2 _6001_/C sky130_fd_sc_hd__a21bo_1
X_4192_ _4303_/A _4192_/B vssd2 vssd2 vccd2 vccd2 _4196_/A sky130_fd_sc_hd__nand2_1
X_6902_ _6834_/A _6834_/B _6832_/X vssd2 vssd2 vccd2 vccd2 _6904_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_77_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7882_ _7886_/CLK _7882_/D _7641_/Y vssd2 vssd2 vccd2 vccd2 _7882_/Q sky130_fd_sc_hd__dfrtp_2
X_6833_ _6833_/A _6833_/B vssd2 vssd2 vccd2 vccd2 _6834_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_525 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_15_92 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7429__S _7451_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6764_ _6694_/A _6612_/Y _6694_/B vssd2 vssd2 vccd2 vccd2 _6767_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_92_539 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3976_ _4454_/A _4018_/A _4018_/B _4164_/C _4328_/A vssd2 vssd2 vccd2 vccd2 _3976_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4042__A1 _4268_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6695_ _6695_/A _6765_/C vssd2 vssd2 vccd2 vccd2 _6769_/C sky130_fd_sc_hd__xor2_1
XANTENNA__6319__B1 _7034_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_72_241 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5715_ _6100_/D _6587_/B _5938_/C vssd2 vssd2 vccd2 vccd2 _5944_/C sky130_fd_sc_hd__and3_2
XFILLER_0_93_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5646_ _7856_/Q _5647_/B vssd2 vssd2 vccd2 vccd2 _5648_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_31_91 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_60_458 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_5_585 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xhold220 hold408/X vssd2 vssd2 vccd2 vccd2 input98/A sky130_fd_sc_hd__dlygate4sd3_1
X_5577_ _7859_/Q _7860_/Q vssd2 vssd2 vccd2 vccd2 _5581_/B sky130_fd_sc_hd__or2_4
XFILLER_0_32_149 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4528_ _4962_/A _4966_/A _4662_/B _4965_/B vssd2 vssd2 vccd2 vccd2 _4529_/B sky130_fd_sc_hd__or4_1
X_7316_ _7316_/A _7316_/B vssd2 vssd2 vccd2 vccd2 _7319_/B sky130_fd_sc_hd__xnor2_1
Xhold253 _7734_/Q vssd2 vssd2 vccd2 vccd2 hold253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 _7736_/Q vssd2 vssd2 vccd2 vccd2 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 _7459_/X vssd2 vssd2 vccd2 vccd2 _7699_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_385 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold286 hold286/A vssd2 vssd2 vccd2 vccd2 la_data_out[26] sky130_fd_sc_hd__buf_12
Xhold275 hold626/X vssd2 vssd2 vccd2 vccd2 hold627/A sky130_fd_sc_hd__dlygate4sd3_1
X_7247_ _7247_/A _7247_/B vssd2 vssd2 vccd2 vccd2 _7279_/B sky130_fd_sc_hd__and2_1
Xhold264 hold264/A vssd2 vssd2 vccd2 vccd2 la_data_out[4] sky130_fd_sc_hd__buf_12
XANTENNA__4089__A _4747_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4459_ _4328_/A _4656_/C _4146_/B _4162_/A vssd2 vssd2 vccd2 vccd2 _4459_/Y sky130_fd_sc_hd__a22oi_1
Xhold297 hold646/X vssd2 vssd2 vccd2 vccd2 hold647/A sky130_fd_sc_hd__dlygate4sd3_1
X_7178_ _7237_/A _7255_/B vssd2 vssd2 vccd2 vccd2 _7179_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_99_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6129_ _6091_/A _6090_/A _6090_/B vssd2 vssd2 vccd2 vccd2 _6142_/A sky130_fd_sc_hd__a21bo_1
XTAP_580 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_149 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_68_569 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_83_528 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_48_282 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_36_433 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_106_321 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_91_572 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_91_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_365 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_63_285 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_51_425 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_23_116 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6479__A _6783_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7038__A1 _7037_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6013__A2 _6664_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_74_539 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5221__B1 _4814_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3830_ _7801_/Q _3831_/B vssd2 vssd2 vccd2 vccd2 _3830_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_109_181 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_82_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_42_403 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5500_ _5500_/A _5500_/B vssd2 vssd2 vccd2 vccd2 _5503_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_488 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6480_ _6707_/A _7181_/A vssd2 vssd2 vccd2 vccd2 _6481_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_42_436 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_14_138 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_499 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_42_469 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_2_500 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5431_ _5431_/A _5431_/B vssd2 vssd2 vccd2 vccd2 _5433_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_112_357 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_2_566 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5362_ _5404_/A _5406_/A _5498_/A _5528_/A vssd2 vssd2 vccd2 vccd2 _5363_/B sky130_fd_sc_hd__or4_1
X_7101_ _7237_/A _7181_/A _7054_/A _7051_/X vssd2 vssd2 vccd2 vccd2 _7103_/B sky130_fd_sc_hd__o31ai_2
X_4313_ _7766_/Q _3982_/B _4032_/C _7769_/Q _4312_/Y vssd2 vssd2 vccd2 vccd2 _4313_/X
+ sky130_fd_sc_hd__a221o_1
X_7032_ _7083_/B _7032_/B vssd2 vssd2 vccd2 vccd2 _7131_/A sky130_fd_sc_hd__or2_2
X_5293_ _5293_/A _5293_/B vssd2 vssd2 vccd2 vccd2 _5293_/Y sky130_fd_sc_hd__xnor2_1
X_4244_ _4244_/A _4299_/A vssd2 vssd2 vccd2 vccd2 _4303_/C sky130_fd_sc_hd__or2_1
X_4175_ _4017_/A _4017_/B _5029_/A vssd2 vssd2 vccd2 vccd2 _4177_/B sky130_fd_sc_hd__a21oi_2
XTAP_1009 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout264_A _7849_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_89_193 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6571__B _6571_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7865_ _7870_/CLK _7865_/D _7624_/Y vssd2 vssd2 vccd2 vccd2 _7865_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_377 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6816_ _6814_/Y _6815_/X _6668_/A _6669_/X vssd2 vssd2 vccd2 vccd2 _6819_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__4015__A1 _7766_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7796_ _7800_/CLK _7796_/D _7555_/Y vssd2 vssd2 vccd2 vccd2 _7796_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__5468__A _5468_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6747_ _6681_/A _6681_/B _6679_/Y vssd2 vssd2 vccd2 vccd2 _6749_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__4015__B2 _7768_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3959_ _4022_/B _4162_/B _4214_/B _4214_/C vssd2 vssd2 vccd2 vccd2 _3967_/C sky130_fd_sc_hd__nor4_1
XFILLER_0_18_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6678_ _6596_/A _6596_/B _6594_/X vssd2 vssd2 vccd2 vccd2 _6680_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_45_296 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_18_488 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5629_ _7862_/Q _5629_/B vssd2 vssd2 vccd2 vccd2 _5664_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_103_357 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_68_300 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1532 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_61 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_72 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1587 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_64_583 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_36_296 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_51_233 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_51_277 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6937__A _6989_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_47_79 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5980_ _6397_/A _5826_/B _5976_/X _5979_/X vssd2 vssd2 vccd2 vccd2 _5980_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_87_653 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_86_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_4931_ _4779_/A _5431_/B _4930_/Y vssd2 vssd2 vccd2 vccd2 _4986_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_63_78 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__5993__A1 _6093_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5993__B2 _6282_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_174 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4862_ _4860_/X _4862_/B vssd2 vssd2 vccd2 vccd2 _4864_/A sky130_fd_sc_hd__and2b_1
X_7650_ _7800_/CLK _7650_/D vssd2 vssd2 vccd2 vccd2 _7650_/Q sky130_fd_sc_hd__dfxtp_1
X_6601_ _6524_/A _6524_/B _6522_/Y vssd2 vssd2 vccd2 vccd2 _6603_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_7_625 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3813_ _3813_/A _3813_/B vssd2 vssd2 vccd2 vccd2 _4457_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_103_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7581_ _7590_/A vssd2 vssd2 vccd2 vccd2 _7581_/Y sky130_fd_sc_hd__inv_2
X_4793_ _4793_/A _4793_/B vssd2 vssd2 vccd2 vccd2 _4830_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_62_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6532_ _6533_/A _6533_/B vssd2 vssd2 vccd2 vccd2 _6610_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_15_436 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6463_ _6392_/A _6392_/B _6318_/A _6317_/B vssd2 vssd2 vccd2 vccd2 _6466_/B sky130_fd_sc_hd__o211ai_1
XFILLER_0_112_121 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5414_ _5414_/A _5414_/B _5528_/A _5528_/B vssd2 vssd2 vccd2 vccd2 _5462_/A sky130_fd_sc_hd__or4_1
Xoutput122 hold657/X vssd2 vssd2 vccd2 vccd2 hold304/A sky130_fd_sc_hd__buf_6
XFILLER_0_112_165 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6394_ _6381_/A _6381_/B _6379_/Y vssd2 vssd2 vccd2 vccd2 _6455_/A sky130_fd_sc_hd__a21oi_2
Xoutput111 hold627/X vssd2 vssd2 vccd2 vccd2 hold276/A sky130_fd_sc_hd__buf_6
XFILLER_0_88_97 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xoutput133 _7646_/Q vssd2 vssd2 vccd2 vccd2 wbs_ack_o sky130_fd_sc_hd__buf_12
XFILLER_0_2_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_56_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5345_ _5297_/A _5296_/B _5294_/X vssd2 vssd2 vccd2 vccd2 _5347_/B sky130_fd_sc_hd__a21oi_1
Xoutput144 _7714_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[19] sky130_fd_sc_hd__buf_12
Xoutput155 _7724_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[29] sky130_fd_sc_hd__buf_12
X_5276_ _5276_/A _5468_/A vssd2 vssd2 vccd2 vccd2 _5279_/A sky130_fd_sc_hd__or2_1
X_7015_ _6961_/A _6960_/B _6960_/A vssd2 vssd2 vccd2 vccd2 _7017_/B sky130_fd_sc_hd__o21ba_1
X_4227_ _4228_/A _4228_/B vssd2 vssd2 vccd2 vccd2 _4227_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_97_406 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4158_ _4229_/A _4229_/B vssd2 vssd2 vccd2 vccd2 _4183_/A sky130_fd_sc_hd__xnor2_1
X_4089_ _4747_/A _4863_/A vssd2 vssd2 vccd2 vccd2 _4090_/C sky130_fd_sc_hd__or2_1
XFILLER_0_77_163 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_92_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7848_ _7854_/CLK _7848_/D _7607_/Y vssd2 vssd2 vccd2 vccd2 _7848_/Q sky130_fd_sc_hd__dfrtp_2
X_7779_ _7779_/CLK _7779_/D _7538_/Y vssd2 vssd2 vccd2 vccd2 _7779_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_92_177 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_73_380 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_46_572 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_61_553 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5645__B _5645_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_61_597 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_21_417 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_33_277 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_33_288 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_21_439 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_108_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_88_417 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5975__A1 _6158_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1340 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_152 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_68_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_33_26 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1384 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_325 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1395 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_177 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5836__A _6670_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xinput13 input13/A vssd2 vssd2 vccd2 vccd2 input13/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_391 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
Xinput35 input35/A vssd2 vssd2 vccd2 vccd2 input35/X sky130_fd_sc_hd__clkbuf_1
Xinput46 input46/A vssd2 vssd2 vccd2 vccd2 input46/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_244 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xinput24 input24/A vssd2 vssd2 vccd2 vccd2 input24/X sky130_fd_sc_hd__clkbuf_1
Xinput57 wbs_adr_i[16] vssd2 vssd2 vccd2 vccd2 _7344_/B sky130_fd_sc_hd__clkbuf_1
Xinput68 input68/A vssd2 vssd2 vccd2 vccd2 input68/X sky130_fd_sc_hd__clkbuf_1
Xinput79 wbs_adr_i[7] vssd2 vssd2 vccd2 vccd2 _7342_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_266 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6089__D _6855_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5130_ _5250_/B _5130_/B vssd2 vssd2 vccd2 vccd2 _5133_/D sky130_fd_sc_hd__xnor2_4
XFILLER_0_20_472 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5061_ _4986_/A _4986_/B _4984_/Y vssd2 vssd2 vccd2 vccd2 _5063_/B sky130_fd_sc_hd__a21oi_2
X_4012_ _4082_/B _4201_/D _4009_/X _4380_/B _7764_/Q vssd2 vssd2 vccd2 vccd2 _4012_/Y
+ sky130_fd_sc_hd__a32oi_1
XFILLER_0_74_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_28_7 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_79_428 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4218__A1 _4598_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5963_ _6059_/A _5963_/B vssd2 vssd2 vccd2 vccd2 _5969_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_87_461 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4914_ _4915_/A _4915_/B vssd2 vssd2 vccd2 vccd2 _4914_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4634__B _4711_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_163 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_59_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7702_ _7782_/CLK _7702_/D vssd2 vssd2 vccd2 vccd2 _7702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_65 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_75_645 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_59_196 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_47_347 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5894_ _6510_/A _5938_/C vssd2 vssd2 vccd2 vccd2 _5894_/X sky130_fd_sc_hd__and2_1
X_4845_ _4845_/A _4845_/B vssd2 vssd2 vccd2 vccd2 _4849_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_7_422 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7633_ _7641_/A vssd2 vssd2 vccd2 vccd2 _7633_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7437__S _7451_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4776_ _5011_/A _5142_/C _5076_/D _4863_/A vssd2 vssd2 vccd2 vccd2 _4778_/A sky130_fd_sc_hd__o22ai_2
X_7564_ _7564_/A vssd2 vssd2 vccd2 vccd2 _7564_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5746__A _7845_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6515_ _6515_/A _6515_/B vssd2 vssd2 vccd2 vccd2 _6516_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout227_A _4880_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_113_441 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7495_ _7524_/A vssd2 vssd2 vccd2 vccd2 _7495_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_255 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6446_ _6446_/A _6446_/B vssd2 vssd2 vccd2 vccd2 _6449_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_236 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_30_247 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_113_485 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6377_ _6377_/A _6377_/B vssd2 vssd2 vccd2 vccd2 _6380_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_461 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5328_ _5328_/A _5528_/B _5458_/C vssd2 vssd2 vccd2 vccd2 _5329_/B sky130_fd_sc_hd__or3_1
XANTENNA__4809__B _4809_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5259_ _5260_/A _5260_/B vssd2 vssd2 vccd2 vccd2 _5349_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__4097__A _5455_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6851__C1 _5781_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_225 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_78_461 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_78_494 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_65_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_93_464 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_66_667 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_19_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_53_328 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_80_158 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_34_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_104_474 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_21_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_21_247 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_409 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
Xfanout190 _4492_/Y vssd2 vssd2 vccd2 vccd2 _5142_/C sky130_fd_sc_hd__clkbuf_8
XANTENNA__4735__A _4966_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_57_623 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_29_314 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1192 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_615 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4630_ _4736_/A _5142_/C _5076_/D _4708_/A vssd2 vssd2 vccd2 vccd2 _4631_/B sky130_fd_sc_hd__o22ai_2
XFILLER_0_44_339 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_114_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5285__B _5550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_114_249 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6300_ _6238_/A _6238_/B _6236_/Y vssd2 vssd2 vccd2 vccd2 _6302_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_80_670 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4561_ _4898_/A _5142_/C vssd2 vssd2 vccd2 vccd2 _4570_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_71_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_52_372 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
Xhold627 hold627/A vssd2 vssd2 vccd2 vccd2 hold627/X sky130_fd_sc_hd__dlygate4sd3_1
X_7280_ _7216_/A _7216_/B _7216_/C _7279_/Y vssd2 vssd2 vccd2 vccd2 _7283_/B sky130_fd_sc_hd__a31o_1
Xhold616 _7811_/Q vssd2 vssd2 vccd2 vccd2 hold616/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold605 hold93/X vssd2 vssd2 vccd2 vccd2 input23/A sky130_fd_sc_hd__dlygate4sd3_1
X_4492_ _4489_/X _4491_/X _4125_/B vssd2 vssd2 vccd2 vccd2 _4492_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_433 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_100_41 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold649 hold649/A vssd2 vssd2 vccd2 vccd2 hold649/X sky130_fd_sc_hd__dlygate4sd3_1
X_6231_ _6233_/A _6233_/B vssd2 vssd2 vccd2 vccd2 _6231_/Y sky130_fd_sc_hd__nand2_1
Xhold638 _7815_/Q vssd2 vssd2 vccd2 vccd2 hold638/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_85 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6162_ _6590_/A _7094_/A vssd2 vssd2 vccd2 vccd2 _6164_/B sky130_fd_sc_hd__nand2_1
XTAP_910 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4629__B _4736_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5113_ _5114_/B _5114_/A vssd2 vssd2 vccd2 vccd2 _5113_/X sky130_fd_sc_hd__and2b_1
XTAP_943 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_291 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_987 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _6093_/A _6152_/B _6152_/C _6102_/B vssd2 vssd2 vccd2 vccd2 _6093_/X sky130_fd_sc_hd__and4_1
XTAP_998 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5044_/A _5044_/B vssd2 vssd2 vccd2 vccd2 _5047_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_79_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_19_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA_fanout177_A _4708_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6995_ _6995_/A _6995_/B vssd2 vssd2 vccd2 vccd2 _6997_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_431 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5946_ _7847_/Q _6281_/B _6281_/C _5853_/B _5853_/C vssd2 vssd2 vccd2 vccd2 _5947_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_464 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_75_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_48_667 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5877_ _6283_/A _5977_/B _5873_/X _5886_/A _5876_/X vssd2 vssd2 vccd2 vccd2 _5883_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_90_401 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_75_486 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4828_ _4829_/B _4829_/A vssd2 vssd2 vccd2 vccd2 _4828_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_62_114 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_47_177 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7616_ _7641_/A vssd2 vssd2 vccd2 vccd2 _7616_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4380__A _4454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_105_205 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_90_467 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_90_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_16_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_16_542 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_28_380 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_105_249 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4759_ _4760_/A _4760_/B vssd2 vssd2 vccd2 vccd2 _4759_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_50_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7547_ _7565_/A vssd2 vssd2 vccd2 vccd2 _7547_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_70_180 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7478_ _7718_/Q _7483_/A2 _7483_/B1 hold343/X vssd2 vssd2 vccd2 vccd2 _7478_/X sky130_fd_sc_hd__a22o_1
X_6429_ _6500_/B _6429_/B vssd2 vssd2 vccd2 vccd2 _6442_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_31_556 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_113_293 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_wb_clk_i clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7806_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5627__B1 _5645_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6570__A1_N _6571_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_98_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__6770__A _7034_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_38_100 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_220 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_109_511 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_54_604 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_38_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_38_155 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_109_555 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_93_261 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_81_423 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_81_401 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_26_328 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_38_166 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_38_188 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_53_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_22_512 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_239 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 hold2/A vssd2 vssd2 vccd2 vccd2 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_501 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6664__B _7099_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_79 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6043__B1 _6150_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6780_ _5994_/X _7222_/A _7222_/C _5948_/X vssd2 vssd2 vccd2 vccd2 _6782_/A sky130_fd_sc_hd__a22o_1
X_3992_ _4598_/A _4747_/A vssd2 vssd2 vccd2 vccd2 _7727_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_29_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5800_ _6158_/A _5977_/B vssd2 vssd2 vccd2 vccd2 _5800_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_57_442 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5731_ _7875_/Q _5731_/B vssd2 vssd2 vccd2 vccd2 _5755_/C sky130_fd_sc_hd__xor2_4
XFILLER_0_29_155 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_29_177 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_29_188 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_72_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_44_136 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5662_ _6093_/A _6194_/B _5662_/C _5662_/D vssd2 vssd2 vccd2 vccd2 _5674_/B sky130_fd_sc_hd__and4_1
X_4613_ _4613_/A _4613_/B vssd2 vssd2 vccd2 vccd2 _4614_/B sky130_fd_sc_hd__xor2_2
X_5593_ _5594_/B _5594_/C vssd2 vssd2 vccd2 vccd2 _6474_/A sky130_fd_sc_hd__and2_2
X_7401_ _7440_/A _7401_/B vssd2 vssd2 vccd2 vccd2 _7669_/D sky130_fd_sc_hd__and2_1
XFILLER_0_111_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7332_ _7335_/A _7325_/Y _7335_/B _7336_/A vssd2 vssd2 vccd2 vccd2 _7333_/B sky130_fd_sc_hd__o31a_1
X_4544_ _4545_/A _4545_/B vssd2 vssd2 vccd2 vccd2 _4618_/A sky130_fd_sc_hd__nand2b_1
Xhold402 hold694/X vssd2 vssd2 vccd2 vccd2 _7802_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_383 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7263_ _7302_/A vssd2 vssd2 vccd2 vccd2 _7263_/Y sky130_fd_sc_hd__inv_2
Xhold424 la_data_in[38] vssd2 vssd2 vccd2 vccd2 hold29/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 hold34/X vssd2 vssd2 vccd2 vccd2 _7844_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 _7869_/Q vssd2 vssd2 vccd2 vccd2 _3804_/A sky130_fd_sc_hd__buf_1
XFILLER_0_40_331 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_96_53 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6214_ _6664_/A _5994_/X _6150_/B _5931_/C vssd2 vssd2 vccd2 vccd2 _6216_/A sky130_fd_sc_hd__a22o_1
X_4475_ _4475_/A _4475_/B vssd2 vssd2 vccd2 vccd2 _4478_/A sky130_fd_sc_hd__xnor2_2
Xhold457 hold15/X vssd2 vssd2 vccd2 vccd2 input28/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 la_data_in[8] vssd2 vssd2 vccd2 vccd2 hold7/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 input4/X vssd2 vssd2 vccd2 vccd2 hold18/A sky130_fd_sc_hd__dlygate4sd3_1
X_7194_ _7140_/A _7255_/B _7141_/A _7139_/B vssd2 vssd2 vccd2 vccd2 _7196_/B sky130_fd_sc_hd__o31a_1
Xhold479 hold14/X vssd2 vssd2 vccd2 vccd2 _7859_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_97 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6145_ _6634_/B _6738_/A vssd2 vssd2 vccd2 vccd2 _6149_/A sky130_fd_sc_hd__nand2_2
XANTENNA__6855__A _6855_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_751 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6093_/A _6194_/C _6130_/C vssd2 vssd2 vccd2 vccd2 _6078_/C sky130_fd_sc_hd__and3_1
X_5027_ _5027_/A _5027_/B vssd2 vssd2 vccd2 vccd2 _5056_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__5085__A1 _5328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_95_515 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_95_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_95_548 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6978_ _6979_/A _6979_/B vssd2 vssd2 vccd2 vccd2 _7060_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_464 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5929_ _5923_/X _5924_/X _5928_/X _5878_/B vssd2 vssd2 vccd2 vccd2 _6425_/A sky130_fd_sc_hd__o31a_4
XFILLER_0_63_434 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_8_572 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_136 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_90_253 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5934__A _6092_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_50_128 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_31_386 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_31_397 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_25_16 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_86_515 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_25_38 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_39_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6328__A1 _6402_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_94_592 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_54_434 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5547__C _5547_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_26_125 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_26_136 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_109_385 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_41_106 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_81_286 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5844__A _6402_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5000__A1 _5133_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5551__A2 _4814_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4260_ _4260_/A _4260_/B _4260_/C vssd2 vssd2 vccd2 vccd2 _4261_/B sky130_fd_sc_hd__nor3_1
XANTENNA__4511__B1 _5222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4191_ _4189_/A _4189_/B _4189_/C _4242_/A _4188_/X vssd2 vssd2 vccd2 vccd2 _4192_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_66_67 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_89_342 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_82_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6901_ _6901_/A _6901_/B vssd2 vssd2 vccd2 vccd2 _6904_/A sky130_fd_sc_hd__xnor2_2
X_7881_ _7886_/CLK _7881_/D _7640_/Y vssd2 vssd2 vccd2 vccd2 _7881_/Q sky130_fd_sc_hd__dfrtp_4
X_6832_ _6833_/A _6833_/B vssd2 vssd2 vccd2 vccd2 _6832_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_99 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_77_537 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_92_507 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4578__B1 _5315_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6763_ _6763_/A _6763_/B vssd2 vssd2 vccd2 vccd2 _7025_/A sky130_fd_sc_hd__xnor2_1
X_3975_ _4125_/C _4021_/D vssd2 vssd2 vccd2 vccd2 _3975_/X sky130_fd_sc_hd__and2_1
X_6694_ _6694_/A _6694_/B vssd2 vssd2 vccd2 vccd2 _6765_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_592 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_9_369 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5714_ _5691_/A _5691_/B _6094_/B vssd2 vssd2 vccd2 vccd2 _5938_/C sky130_fd_sc_hd__a21oi_4
XFILLER_0_5_520 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5645_ _7855_/Q _5645_/B vssd2 vssd2 vccd2 vccd2 _5647_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_33_607 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_86_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_60_415 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7445__S _7451_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_13_320 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold210 _7425_/X vssd2 vssd2 vccd2 vccd2 _7426_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5576_ _7856_/Q _7855_/Q _7857_/Q _7858_/Q vssd2 vssd2 vccd2 vccd2 _5581_/A sky130_fd_sc_hd__or4_4
XANTENNA__6288__C _6430_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4527_ _4966_/A _4662_/B _4965_/B _4962_/A vssd2 vssd2 vccd2 vccd2 _4527_/X sky130_fd_sc_hd__o22a_1
X_7315_ _7315_/A _7315_/B vssd2 vssd2 vccd2 vccd2 _7316_/B sky130_fd_sc_hd__nor2_1
Xhold221 input98/X vssd2 vssd2 vccd2 vccd2 hold221/X sky130_fd_sc_hd__buf_1
Xhold232 _7464_/X vssd2 vssd2 vccd2 vccd2 _7704_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 _7735_/Q vssd2 vssd2 vccd2 vccd2 hold243/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold276 hold276/A vssd2 vssd2 vccd2 vccd2 la_data_out[19] sky130_fd_sc_hd__buf_12
Xhold287 hold638/X vssd2 vssd2 vccd2 vccd2 hold639/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 hold618/X vssd2 vssd2 vccd2 vccd2 hold619/A sky130_fd_sc_hd__dlygate4sd3_1
X_7246_ _7246_/A _7246_/B _7246_/C vssd2 vssd2 vccd2 vccd2 _7247_/B sky130_fd_sc_hd__or3_1
Xhold254 _7462_/X vssd2 vssd2 vccd2 vccd2 _7702_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4089__B _4863_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4458_ _4814_/A _4519_/B _4458_/C _4458_/D vssd2 vssd2 vccd2 vccd2 _4458_/X sky130_fd_sc_hd__or4_1
Xhold298 hold298/A vssd2 vssd2 vccd2 vccd2 la_data_out[15] sky130_fd_sc_hd__buf_12
XANTENNA__6585__A _6668_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7177_ _7177_/A _7177_/B vssd2 vssd2 vccd2 vccd2 _7179_/A sky130_fd_sc_hd__nand2_1
X_6128_ _6128_/A _6128_/B _6128_/C vssd2 vssd2 vccd2 vccd2 _6182_/A sky130_fd_sc_hd__and3_1
X_4389_ _4962_/A _5042_/A _4662_/B _5042_/B vssd2 vssd2 vccd2 vccd2 _4390_/B sky130_fd_sc_hd__or4_1
XTAP_570 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _6059_/A _6064_/B _6128_/A _6059_/D vssd2 vssd2 vccd2 vccd2 _6062_/A sky130_fd_sc_hd__nor4_2
XFILLER_0_95_345 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_68_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_48_261 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_36_401 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_36_412 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_48_294 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_11_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_333 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_91_584 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_51_437 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7355__S _7383_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5664__A _6157_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_106_377 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6479__B _6855_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_32_662 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6495__A _6989_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7038__A2 _7253_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_99_662 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_86_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5839__A _6093_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_356 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_59_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_74_529 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_27_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_54_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_109_193 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_54_275 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5430_ _5430_/A _5430_/B vssd2 vssd2 vccd2 vccd2 _5433_/B sky130_fd_sc_hd__xnor2_1
X_5361_ _5081_/C _5498_/A _5528_/A _5404_/A vssd2 vssd2 vccd2 vccd2 _5363_/A sky130_fd_sc_hd__o22ai_1
X_7100_ _7100_/A _7100_/B vssd2 vssd2 vccd2 vccd2 _7103_/A sky130_fd_sc_hd__xnor2_1
X_5292_ _5292_/A _5292_/B vssd2 vssd2 vccd2 vccd2 _5293_/B sky130_fd_sc_hd__xnor2_2
X_4312_ _4312_/A _4814_/B vssd2 vssd2 vccd2 vccd2 _4312_/Y sky130_fd_sc_hd__nor2_1
X_7031_ _7211_/A _7031_/B _7031_/C vssd2 vssd2 vccd2 vccd2 _7032_/B sky130_fd_sc_hd__and3_1
X_4243_ _4243_/A _4243_/B vssd2 vssd2 vccd2 vccd2 _4299_/A sky130_fd_sc_hd__nor2_1
X_4174_ _4044_/A _4044_/B _5042_/A vssd2 vssd2 vccd2 vccd2 _4177_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_109 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_89_161 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA_fanout257_A _7853_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7864_ _7870_/CLK _7864_/D _7623_/Y vssd2 vssd2 vccd2 vccd2 _7864_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_58_570 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6815_ _6815_/A _6815_/B _6815_/C vssd2 vssd2 vccd2 vccd2 _6815_/X sky130_fd_sc_hd__and3_1
X_7795_ _7795_/CLK _7795_/D _7554_/Y vssd2 vssd2 vccd2 vccd2 _7795_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5468__B _5550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6746_ _6746_/A _6746_/B vssd2 vssd2 vccd2 vccd2 _6749_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_220 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_73_540 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_9_177 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_18_467 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3958_ _4162_/B _4214_/B vssd2 vssd2 vccd2 vccd2 _3986_/A sky130_fd_sc_hd__nor2_1
X_6677_ _6677_/A _6677_/B vssd2 vssd2 vccd2 vccd2 _6680_/A sky130_fd_sc_hd__xnor2_2
X_3889_ _7792_/Q _3889_/B vssd2 vssd2 vccd2 vccd2 _3893_/D sky130_fd_sc_hd__xor2_2
X_5628_ _7862_/Q _5629_/B vssd2 vssd2 vccd2 vccd2 _6019_/C sky130_fd_sc_hd__xor2_4
X_5559_ _5570_/A _5559_/B vssd2 vssd2 vccd2 vccd2 _5573_/C sky130_fd_sc_hd__or2_1
XANTENNA__6476__B1 _7222_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5931__B _6402_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_111_391 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7229_ _7229_/A _7229_/B vssd2 vssd2 vccd2 vccd2 _7230_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_96_610 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1533 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_507 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_62 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_73 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_337 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_95 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_84 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_106_141 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_36_264 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_51_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_24_448 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_20_610 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6937__B _7253_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_47_36 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__6219__B1 _7045_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_78_109 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_99_470 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_63_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_87_665 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4930_ _4930_/A _4930_/B vssd2 vssd2 vccd2 vccd2 _4930_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_345 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_87_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4861_ _5042_/A _5168_/A _5142_/C _5076_/D vssd2 vssd2 vccd2 vccd2 _4862_/B sky130_fd_sc_hd__or4_1
XFILLER_0_59_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6600_ _6600_/A _6600_/B vssd2 vssd2 vccd2 vccd2 _6603_/A sky130_fd_sc_hd__xnor2_2
X_3812_ _3813_/A _3813_/B vssd2 vssd2 vccd2 vccd2 _4519_/B sky130_fd_sc_hd__and2_4
X_7580_ _7590_/A vssd2 vssd2 vccd2 vccd2 _7580_/Y sky130_fd_sc_hd__inv_2
X_4792_ _4793_/B _4793_/A vssd2 vssd2 vccd2 vccd2 _4854_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_7_648 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6531_ _6531_/A _6531_/B vssd2 vssd2 vccd2 vccd2 _6533_/B sky130_fd_sc_hd__xor2_2
XANTENNA__4953__B1 _5550_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_6_136 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6462_ _6615_/A _6462_/B vssd2 vssd2 vccd2 vccd2 _6466_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_42_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_112_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6393_ _6393_/A _6393_/B vssd2 vssd2 vccd2 vccd2 _7818_/D sky130_fd_sc_hd__xnor2_1
Xoutput101 hold609/X vssd2 vssd2 vccd2 vccd2 hold256/A sky130_fd_sc_hd__buf_6
XFILLER_0_70_587 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_42_278 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5413_ _5326_/B _5030_/C _4814_/Y _4800_/C vssd2 vssd2 vccd2 vccd2 _5415_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_88_65 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xoutput123 hold623/X vssd2 vssd2 vccd2 vccd2 hold270/A sky130_fd_sc_hd__buf_6
Xoutput112 hold615/X vssd2 vssd2 vccd2 vccd2 hold262/A sky130_fd_sc_hd__buf_6
X_5344_ _5344_/A _5344_/B vssd2 vssd2 vccd2 vccd2 _5347_/A sky130_fd_sc_hd__xnor2_1
Xoutput134 _7695_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[0] sky130_fd_sc_hd__buf_12
XFILLER_0_112_177 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_11_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xoutput145 _7696_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[1] sky130_fd_sc_hd__buf_12
Xoutput156 _7697_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[2] sky130_fd_sc_hd__buf_12
X_5275_ _5275_/A _5275_/B vssd2 vssd2 vccd2 vccd2 _5293_/A sky130_fd_sc_hd__xor2_2
XANTENNA__7024__A _7024_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7014_ _7014_/A _7014_/B vssd2 vssd2 vccd2 vccd2 _7017_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4226_ _4226_/A _4226_/B vssd2 vssd2 vccd2 vccd2 _4228_/B sky130_fd_sc_hd__xnor2_1
X_4157_ _4229_/A _4229_/B vssd2 vssd2 vccd2 vccd2 _4230_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_69_109 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4088_ _4088_/A _4088_/B vssd2 vssd2 vccd2 vccd2 _4736_/A sky130_fd_sc_hd__and2_2
XFILLER_0_78_654 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4383__A _7770_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_93_613 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_77_153 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7847_ _7854_/CLK _7847_/D _7606_/Y vssd2 vssd2 vccd2 vccd2 _7847_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5198__B _5357_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_80_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_46_562 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7778_ _7779_/CLK _7778_/D _7537_/Y vssd2 vssd2 vccd2 vccd2 _7778_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_220 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_92_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6729_ _6729_/A _6729_/B vssd2 vssd2 vccd2 vccd2 _6731_/A sky130_fd_sc_hd__nand2_1
Xwire239 _4020_/B vssd2 vssd2 vccd2 vccd2 _4125_/C sky130_fd_sc_hd__buf_2
Xwire228 _3902_/Y vssd2 vssd2 vccd2 vccd2 wire228/X sky130_fd_sc_hd__buf_1
XFILLER_0_103_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_61_565 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_14_481 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5942__A _6093_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_17_28 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_88_429 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6621__B1 _7034_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4576__C_N _5030_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1341 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_518 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_38 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1374 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_197 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_68_186 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XTAP_1396 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_107_472 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6137__C1 _5736_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xinput36 input36/A vssd2 vssd2 vccd2 vccd2 input36/X sky130_fd_sc_hd__clkbuf_1
Xinput25 input25/A vssd2 vssd2 vccd2 vccd2 input25/X sky130_fd_sc_hd__clkbuf_1
Xinput14 input14/A vssd2 vssd2 vccd2 vccd2 input14/X sky130_fd_sc_hd__buf_1
XFILLER_0_52_587 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xinput58 wbs_adr_i[17] vssd2 vssd2 vccd2 vccd2 _7344_/A sky130_fd_sc_hd__clkbuf_1
Xinput47 input47/A vssd2 vssd2 vccd2 vccd2 input47/X sky130_fd_sc_hd__clkbuf_1
Xinput69 wbs_adr_i[27] vssd2 vssd2 vccd2 vccd2 _7339_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__5852__A _6253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5360__B1 _5455_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_58_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7101__A1 _7237_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5060_ _5060_/A _5060_/B vssd2 vssd2 vccd2 vccd2 _5063_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_20_495 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4011_ _7767_/Q _4326_/B _4326_/C _4268_/D vssd2 vssd2 vccd2 vccd2 _4011_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_74_45 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5962_ _5962_/A _5962_/B _5962_/C vssd2 vssd2 vccd2 vccd2 _5963_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_59_120 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_87_473 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4913_ _4830_/A _4830_/B _4828_/X vssd2 vssd2 vccd2 vccd2 _4915_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__4634__C _5042_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7701_ _7798_/CLK _7701_/D vssd2 vssd2 vccd2 vccd2 _7701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_87_484 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5893_ _6402_/A _6150_/A vssd2 vssd2 vccd2 vccd2 _5910_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4844_ _4687_/Y _4691_/B _4768_/B _4843_/X vssd2 vssd2 vccd2 vccd2 _4845_/B sky130_fd_sc_hd__o31ai_4
X_7632_ _7641_/A vssd2 vssd2 vccd2 vccd2 _7632_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_412 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_74_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4775_ _4733_/A _4733_/B _4731_/Y vssd2 vssd2 vccd2 vccd2 _4791_/A sky130_fd_sc_hd__a21o_2
XANTENNA__4650__B _4965_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_7_434 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5746__B _6152_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7563_ _7563_/A vssd2 vssd2 vccd2 vccd2 _7563_/Y sky130_fd_sc_hd__inv_2
X_6514_ _6590_/A _6515_/A _7294_/C vssd2 vssd2 vccd2 vccd2 _6514_/X sky130_fd_sc_hd__and3_1
XFILLER_0_43_554 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_43_532 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_70_340 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7494_ _7524_/A vssd2 vssd2 vccd2 vccd2 _7494_/Y sky130_fd_sc_hd__inv_2
X_6445_ _6445_/A _6445_/B vssd2 vssd2 vccd2 vccd2 _6446_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_604 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_70_384 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_3_673 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_113_497 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6376_ _6376_/A _6376_/B vssd2 vssd2 vccd2 vccd2 _6377_/B sky130_fd_sc_hd__xnor2_2
X_5327_ _4965_/B _5528_/B _5458_/C vssd2 vssd2 vccd2 vccd2 _5329_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__4528__D _4965_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5258_ _5206_/A _5208_/B _5206_/B vssd2 vssd2 vccd2 vccd2 _5260_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__6851__B1 _7222_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5189_ _5191_/A _5191_/B vssd2 vssd2 vccd2 vccd2 _5189_/Y sky130_fd_sc_hd__nor2_1
X_4209_ _4807_/A _5042_/A vssd2 vssd2 vccd2 vccd2 _4219_/B sky130_fd_sc_hd__or2_1
XFILLER_0_97_237 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5937__A _6157_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_65_134 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_19_540 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_93_476 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_81_627 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_80_104 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_65_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_65_178 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_148 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_137 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_46_392 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__7363__S _7383_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5342__B1 _5207_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_28_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6842__B1 _7034_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7599__A _7627_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3920__A _7763_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout191 _5366_/A vssd2 vssd2 vccd2 vccd2 _5276_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__4735__B _5220_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_56_123 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XTAP_1182 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_359 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XTAP_1193 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_318 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_37_370 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4560_ _4517_/A _4517_/B _4515_/Y vssd2 vssd2 vccd2 vccd2 _4572_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__4384__A1 _4328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_107_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_4_448 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xhold617 hold617/A vssd2 vssd2 vccd2 vccd2 hold617/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_395 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_12_237 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xhold606 input23/X vssd2 vssd2 vccd2 vccd2 hold94/A sky130_fd_sc_hd__dlygate4sd3_1
X_4491_ _4893_/A _4020_/B _4030_/X _4706_/A1 _4490_/Y vssd2 vssd2 vccd2 vccd2 _4491_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_401 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_100_53 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold628 _7817_/Q vssd2 vssd2 vccd2 vccd2 hold628/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 hold639/A vssd2 vssd2 vccd2 vccd2 hold639/X sky130_fd_sc_hd__dlygate4sd3_1
X_6230_ _6668_/A _6150_/B _6165_/B _6163_/X vssd2 vssd2 vccd2 vccd2 _6233_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_69_78 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_100_97 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_900 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4198__A _4454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6161_ _6152_/X _6153_/X _6159_/X _5944_/B vssd2 vssd2 vccd2 vccd2 _6986_/A sky130_fd_sc_hd__o31ai_4
XANTENNA__7086__B1 _7034_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4629__C _5142_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5112_ _5038_/Y _5052_/B _5050_/Y vssd2 vssd2 vccd2 vccd2 _5114_/B sky130_fd_sc_hd__a21oi_2
XTAP_944 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_85_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6092_ _6092_/A _6939_/A vssd2 vssd2 vccd2 vccd2 _6106_/A sky130_fd_sc_hd__nor2_1
XTAP_977 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XTAP_999 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5041_/X _5043_/B vssd2 vssd2 vccd2 vccd2 _5044_/B sky130_fd_sc_hd__and2b_1
X_6994_ _6995_/A _6995_/B vssd2 vssd2 vccd2 vccd2 _6994_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_87_281 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5945_ _6283_/A _5769_/X _5785_/X _6158_/A _5944_/X vssd2 vssd2 vccd2 vccd2 _5945_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_75_443 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5876_ _7843_/Q _5588_/Y _6398_/B _7844_/Q vssd2 vssd2 vccd2 vccd2 _5876_/X sky130_fd_sc_hd__a22o_1
X_4827_ _4753_/A _4753_/B _4751_/X vssd2 vssd2 vccd2 vccd2 _4829_/B sky130_fd_sc_hd__o21ba_2
XFILLER_0_47_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_16_510 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7615_ _7641_/A vssd2 vssd2 vccd2 vccd2 _7615_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_105_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4375__A1 _4454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4758_ _4677_/A _4677_/B _4675_/X vssd2 vssd2 vccd2 vccd2 _4760_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_80 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7546_ _7563_/A vssd2 vssd2 vccd2 vccd2 _7546_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_286 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6588__A _6670_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7477_ _7717_/Q _7483_/A2 _7483_/B1 hold341/X vssd2 vssd2 vccd2 vccd2 _7477_/X sky130_fd_sc_hd__a22o_1
X_4689_ _4479_/A _4480_/A _4479_/B _4551_/A _4619_/C vssd2 vssd2 vccd2 vccd2 _4689_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_113_261 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_101_401 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6428_ _6738_/A _6571_/C _6427_/C vssd2 vssd2 vccd2 vccd2 _6429_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__4127__B2 _7764_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4127__A1 _7763_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_101_434 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_11_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6100__B _6281_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6359_ _6253_/A _6281_/C _5751_/Y _6093_/A _6358_/Y vssd2 vssd2 vccd2 vccd2 _6359_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_98_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_98_579 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_14_18 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XPHY_210 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_78_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_66_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_14_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_221 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_93_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_54_649 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_30_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_22_524 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_192 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5833__C _6424_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_22_579 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_37 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6945__B _7181_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4746__A _4810_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold3 hold3/A vssd2 vssd2 vccd2 vccd2 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6291__A1 _6668_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_89_557 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_89_568 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_57_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3991_ hold411/X _3981_/X _3990_/X vssd2 vssd2 vccd2 vccd2 _3991_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_9_529 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5730_ _7874_/Q _5730_/B vssd2 vssd2 vccd2 vccd2 _5755_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_29_134 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_57_465 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7400_ hold169/X _7781_/D _7418_/S vssd2 vssd2 vccd2 vccd2 _7400_/X sky130_fd_sc_hd__mux2_1
X_5661_ _7855_/Q _5661_/B _5836_/B _5665_/B vssd2 vssd2 vccd2 vccd2 _5662_/D sky130_fd_sc_hd__and4_1
XFILLER_0_72_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_60_608 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4612_ _4613_/A _4613_/B vssd2 vssd2 vccd2 vccd2 _4612_/Y sky130_fd_sc_hd__nor2_1
X_5592_ _7868_/Q _5598_/B _5592_/C vssd2 vssd2 vccd2 vccd2 _5594_/C sky130_fd_sc_hd__or3_2
X_7331_ _7334_/A _7334_/B _7334_/D vssd2 vssd2 vccd2 vccd2 _7333_/A sky130_fd_sc_hd__and3_1
X_4543_ _4543_/A _4543_/B vssd2 vssd2 vccd2 vccd2 _4545_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_20_50 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_209 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold414 _7337_/X vssd2 vssd2 vccd2 vccd2 _7837_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 la_data_in[43] vssd2 vssd2 vccd2 vccd2 hold31/A sky130_fd_sc_hd__dlygate4sd3_1
X_7262_ _7264_/A _7264_/B vssd2 vssd2 vccd2 vccd2 _7302_/A sky130_fd_sc_hd__nor2_1
Xhold425 hold29/X vssd2 vssd2 vccd2 vccd2 input32/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold403 _7790_/Q vssd2 vssd2 vccd2 vccd2 _4049_/B sky130_fd_sc_hd__buf_1
XANTENNA__5743__C _6670_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_20_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6213_ _6855_/A _6581_/A vssd2 vssd2 vccd2 vccd2 _6217_/A sky130_fd_sc_hd__nor2_1
Xmax_cap166 _6062_/A vssd2 vssd2 vccd2 vccd2 _6122_/B sky130_fd_sc_hd__buf_1
X_4474_ _4474_/A _4474_/B vssd2 vssd2 vccd2 vccd2 _4475_/B sky130_fd_sc_hd__xnor2_2
Xhold469 hold7/X vssd2 vssd2 vccd2 vccd2 input47/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 hold18/X vssd2 vssd2 vccd2 vccd2 _7883_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 input28/X vssd2 vssd2 vccd2 vccd2 hold16/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_253 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_96_65 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7193_ _7153_/A _7191_/B _7151_/Y _7154_/Y vssd2 vssd2 vccd2 vccd2 _7196_/A sky130_fd_sc_hd__o31a_1
XANTENNA__3868__B1 _7764_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6144_ _6144_/A _6144_/B vssd2 vssd2 vccd2 vccd2 _6173_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__6855__B _7255_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_752 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4656__A _4656_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6075_ _6398_/A _6253_/C _6075_/C _6075_/D vssd2 vssd2 vccd2 vccd2 _6078_/B sky130_fd_sc_hd__and4_1
X_5026_ _5027_/B _5027_/A vssd2 vssd2 vccd2 vccd2 _5072_/B sky130_fd_sc_hd__and2b_1
XANTENNA__5085__A2 _5366_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_796 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout287_A _7629_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_31_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_95_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_67_207 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_45_91 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6034__A1 _6282_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6977_ _6977_/A _6977_/B vssd2 vssd2 vccd2 vccd2 _6979_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__6034__B2 _6157_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4045__B1 _4882_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5928_ _6670_/A _5878_/C _5925_/X _5926_/X _5927_/X vssd2 vssd2 vccd2 vccd2 _5928_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_90_221 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_63_446 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5859_ _6158_/A _5769_/X _5785_/X _7847_/Q vssd2 vssd2 vccd2 vccd2 _5859_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_35_126 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_548 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_90_265 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_63_457 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_148 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5934__B _6138_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7529_ _7561_/A vssd2 vssd2 vccd2 vccd2 _7529_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4520__B2 _4809_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4520__A1 _4162_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7470__B1 _7483_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_98_321 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_98_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_98_354 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__6781__A _6855_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_58_229 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_94_571 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6328__A2 _6404_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_54_446 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4339__A1 _4882_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_26_159 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_34_192 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_10_538 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4190_ _4190_/A vssd2 vssd2 vccd2 vccd2 _4303_/A sky130_fd_sc_hd__inv_2
XFILLER_0_66_46 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7461__B1 _7485_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_89_354 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_77_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6900_ _6900_/A _6900_/B vssd2 vssd2 vccd2 vccd2 _6901_/B sky130_fd_sc_hd__xnor2_2
X_7880_ _7886_/CLK _7880_/D _7639_/Y vssd2 vssd2 vccd2 vccd2 _7880_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_106_41 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6831_ _6754_/A _6754_/B _6752_/Y vssd2 vssd2 vccd2 vccd2 _6833_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_82_89 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_49_229 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_85 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6762_ _6762_/A _6762_/B vssd2 vssd2 vccd2 vccd2 _6768_/A sky130_fd_sc_hd__and2_1
XFILLER_0_85_571 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_3974_ _4125_/B _4022_/B _4162_/B _4214_/B vssd2 vssd2 vccd2 vccd2 _4021_/D sky130_fd_sc_hd__nor4_1
X_6693_ _6693_/A _6693_/B vssd2 vssd2 vccd2 vccd2 _6694_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_72_221 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5713_ _6100_/D _6587_/B vssd2 vssd2 vccd2 vccd2 _5713_/Y sky130_fd_sc_hd__nand2_2
X_5644_ _7857_/Q _5644_/B vssd2 vssd2 vccd2 vccd2 _5665_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_72_298 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_5_565 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_32_129 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_79_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7314_ _7253_/C _7291_/B _6670_/Y _7253_/B _7313_/Y vssd2 vssd2 vccd2 vccd2 _7315_/B
+ sky130_fd_sc_hd__o221a_1
Xhold200 hold381/X vssd2 vssd2 vccd2 vccd2 _7779_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 wbs_dat_i[14] vssd2 vssd2 vccd2 vccd2 input88/A sky130_fd_sc_hd__dlygate4sd3_1
X_5575_ _4893_/A _4006_/B hold676/X _7758_/D vssd2 vssd2 vccd2 vccd2 _7757_/D sky130_fd_sc_hd__a31o_1
X_4526_ _4810_/A _5315_/B vssd2 vssd2 vccd2 vccd2 _4530_/A sky130_fd_sc_hd__or2_1
Xhold233 _7739_/Q vssd2 vssd2 vccd2 vccd2 hold233/X sky130_fd_sc_hd__buf_1
Xhold244 _7463_/X vssd2 vssd2 vccd2 vccd2 _7703_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 _7439_/X vssd2 vssd2 vccd2 vccd2 _7440_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout202_A _4217_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_111_573 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xhold277 hold628/X vssd2 vssd2 vccd2 vccd2 hold629/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 hold266/A vssd2 vssd2 vccd2 vccd2 la_data_out[5] sky130_fd_sc_hd__buf_12
Xhold255 hold608/X vssd2 vssd2 vccd2 vccd2 hold609/A sky130_fd_sc_hd__dlygate4sd3_1
X_7245_ _7246_/A _7246_/B _7246_/C vssd2 vssd2 vccd2 vccd2 _7247_/A sky130_fd_sc_hd__o21ai_2
X_4457_ _4457_/A _4457_/B _4458_/C vssd2 vssd2 vccd2 vccd2 _4457_/X sky130_fd_sc_hd__or3_1
Xhold299 hold652/X vssd2 vssd2 vccd2 vccd2 hold653/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 hold288/A vssd2 vssd2 vccd2 vccd2 la_data_out[8] sky130_fd_sc_hd__buf_12
X_7176_ _7224_/A _7253_/A _7291_/A _7253_/B vssd2 vssd2 vccd2 vccd2 _7177_/B sky130_fd_sc_hd__or4_1
X_6127_ _6127_/A _6189_/B vssd2 vssd2 vccd2 vccd2 _7814_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__6585__B _7222_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4388_ _5042_/A _4662_/B _5042_/B _4962_/A vssd2 vssd2 vccd2 vccd2 _4388_/X sky130_fd_sc_hd__o22a_1
XTAP_560 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _6057_/B _6057_/C _6057_/A vssd2 vssd2 vccd2 vccd2 _6059_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__4266__B1 _5458_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5009_ _5168_/A _5207_/A _5142_/C _5076_/D vssd2 vssd2 vccd2 vccd2 _5010_/B sky130_fd_sc_hd__or4_1
XFILLER_0_95_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_95_368 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_48_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_106_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_106_345 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_23_107 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_106_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6479__C _6479_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_16_192 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7371__S _7383_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6495__B _6973_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_86_313 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_59_516 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_52_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_98_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_86_368 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_67_571 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6016__A _7849_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_6_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_109_161 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_54_287 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_42_416 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_42_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_50_471 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5360_ _5454_/A _5454_/B _5455_/A vssd2 vssd2 vccd2 vccd2 _5402_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_2_557 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_77_23 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_50_493 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5291_ _5292_/A _5292_/B vssd2 vssd2 vccd2 vccd2 _5341_/C sky130_fd_sc_hd__and2b_1
XFILLER_0_10_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_22_173 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4311_ _4706_/A1 _4162_/B _4057_/C _7771_/Q _4125_/B vssd2 vssd2 vccd2 vccd2 _4311_/X
+ sky130_fd_sc_hd__a32o_1
X_7030_ _7031_/B _7031_/C _7211_/A vssd2 vssd2 vccd2 vccd2 _7083_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_368 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4242_ _4242_/A _4243_/B vssd2 vssd2 vccd2 vccd2 _4301_/A sky130_fd_sc_hd__or2_1
XANTENNA__5590__A _5645_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4173_ _4598_/A _4729_/A _5030_/B vssd2 vssd2 vccd2 vccd2 _4178_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_93_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5996__B1 _5994_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4934__A _5042_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_26_82 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_26_93 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_77_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6571__D _7094_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7863_ _7870_/CLK _7863_/D _7622_/Y vssd2 vssd2 vccd2 vccd2 _7863_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_65_519 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6814_ _6815_/A _6815_/B _6815_/C vssd2 vssd2 vccd2 vccd2 _6814_/Y sky130_fd_sc_hd__a21oi_1
X_7794_ _7795_/CLK _7794_/D _7553_/Y vssd2 vssd2 vccd2 vccd2 _7794_/Q sky130_fd_sc_hd__dfrtp_4
X_6745_ _6745_/A _6745_/B vssd2 vssd2 vccd2 vccd2 _6746_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_593 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_58_582 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_45_210 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3957_ _4164_/C _5030_/A vssd2 vssd2 vccd2 vccd2 _4018_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_18_413 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6676_ _6676_/A _6676_/B vssd2 vssd2 vccd2 vccd2 _6677_/B sky130_fd_sc_hd__xor2_2
X_3888_ _7791_/Q _3888_/B vssd2 vssd2 vccd2 vccd2 _3889_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_246 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5627_ _7861_/Q _5581_/A _5581_/B _5645_/B vssd2 vssd2 vccd2 vccd2 _5629_/B sky130_fd_sc_hd__o31a_4
XFILLER_0_103_337 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5558_ _5558_/A _5558_/B vssd2 vssd2 vccd2 vccd2 _5559_/B sky130_fd_sc_hd__and2_1
X_4509_ _4729_/A _5042_/B _5030_/B vssd2 vssd2 vccd2 vccd2 _4514_/A sky130_fd_sc_hd__or3b_2
XFILLER_0_13_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_41_482 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_41_493 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6476__A1 _6402_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6476__B2 _5819_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5931__C _5931_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7228_ _7229_/A _7229_/B vssd2 vssd2 vccd2 vccd2 _7259_/B sky130_fd_sc_hd__or2_1
X_5489_ _5488_/A _5488_/B _5518_/B vssd2 vssd2 vccd2 vccd2 _5490_/B sky130_fd_sc_hd__a21oi_1
X_7159_ _7107_/A _7107_/B _7105_/Y vssd2 vssd2 vccd2 vccd2 _7162_/A sky130_fd_sc_hd__a21oi_1
XTAP_390 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_600 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_68_313 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1512 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_52 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_63 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_74 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_349 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_96 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_64_541 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_36_232 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_51_213 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_24_427 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_107_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_106_153 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_91_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_106_197 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_51_257 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_32_471 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_7_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7878_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_47_15 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__6219__A1 _5816_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4860_ _5168_/A _5404_/A _5076_/D _4704_/B vssd2 vssd2 vccd2 vccd2 _4860_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_74_305 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3811_ _7802_/Q _3831_/B _3811_/C vssd2 vssd2 vccd2 vccd2 _3813_/B sky130_fd_sc_hd__or3_4
X_6530_ _6531_/A _6531_/B vssd2 vssd2 vccd2 vccd2 _6610_/A sky130_fd_sc_hd__or2_1
X_4791_ _4791_/A _4791_/B vssd2 vssd2 vccd2 vccd2 _4793_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_67_390 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_55_552 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5585__A _5645_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_27_221 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4953__A1 _5029_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4953__B2 _4882_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6461_ _6461_/A _6461_/B vssd2 vssd2 vccd2 vccd2 _6462_/B sky130_fd_sc_hd__and2_1
XFILLER_0_70_544 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_70_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_15_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_27_298 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6392_ _6392_/A _6392_/B vssd2 vssd2 vccd2 vccd2 _6393_/B sky130_fd_sc_hd__or2_1
XFILLER_0_30_408 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_30_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5412_ _5412_/A _5412_/B vssd2 vssd2 vccd2 vccd2 _5420_/B sky130_fd_sc_hd__nand2_1
Xoutput124 hold633/X vssd2 vssd2 vccd2 vccd2 hold272/A sky130_fd_sc_hd__buf_6
Xoutput113 hold645/X vssd2 vssd2 vccd2 vccd2 hold294/A sky130_fd_sc_hd__buf_6
XFILLER_0_100_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xoutput102 hold629/X vssd2 vssd2 vccd2 vccd2 hold278/A sky130_fd_sc_hd__buf_6
XFILLER_0_88_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5343_ _5344_/B vssd2 vssd2 vccd2 vccd2 _5343_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_112_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
Xoutput135 _7705_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[10] sky130_fd_sc_hd__buf_12
Xoutput146 _7715_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[20] sky130_fd_sc_hd__buf_12
Xoutput157 _7725_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[30] sky130_fd_sc_hd__buf_12
X_5274_ _5275_/A _5275_/B vssd2 vssd2 vccd2 vccd2 _5274_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__7024__B _7024_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7013_ _7012_/A _7012_/B _7012_/C vssd2 vssd2 vccd2 vccd2 _7014_/B sky130_fd_sc_hd__o21ai_1
X_4225_ _4044_/A _4044_/B _4896_/A vssd2 vssd2 vccd2 vccd2 _4226_/B sky130_fd_sc_hd__a21oi_1
X_4156_ _4747_/A _4896_/A vssd2 vssd2 vccd2 vccd2 _4229_/B sky130_fd_sc_hd__nor2_1
XANTENNA__6630__A1 _5819_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4087_ _4081_/X _4082_/X _4087_/C _4087_/D vssd2 vssd2 vccd2 vccd2 _4088_/B sky130_fd_sc_hd__and4bb_2
XFILLER_0_77_110 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4894__A1_N _4810_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7846_ _7854_/CLK _7846_/D _7605_/Y vssd2 vssd2 vccd2 vccd2 _7846_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_647 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_77_187 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4989_ _4989_/A _4989_/B vssd2 vssd2 vccd2 vccd2 _4990_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_46_541 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7777_ _7779_/CLK _7777_/D _7536_/Y vssd2 vssd2 vccd2 vccd2 _7777_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_243 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4944__A1 _5145_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6728_ _6973_/A _6973_/B _7140_/A _7237_/A vssd2 vssd2 vccd2 vccd2 _6729_/B sky130_fd_sc_hd__or4_1
XFILLER_0_18_287 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_104_602 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6146__B1 _5994_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6659_ _6660_/A _6660_/B vssd2 vssd2 vccd2 vccd2 _6659_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_73_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_213 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_235 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_246 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_577 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_14_460 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5942__B _5992_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_103_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_96_463 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1331 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_165 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_68_132 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1375 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_102 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1397 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_658 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_71_319 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_71_308 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6137__B1 _6973_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xinput37 input37/A vssd2 vssd2 vccd2 vccd2 input37/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xinput26 input26/A vssd2 vssd2 vccd2 vccd2 input26/X sky130_fd_sc_hd__clkbuf_1
Xinput15 input15/A vssd2 vssd2 vccd2 vccd2 input15/X sky130_fd_sc_hd__clkbuf_1
Xinput48 input48/A vssd2 vssd2 vccd2 vccd2 input48/X sky130_fd_sc_hd__buf_1
Xinput59 wbs_adr_i[18] vssd2 vssd2 vccd2 vccd2 _7344_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5360__A1 _5454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_58_69 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7101__A2 _7181_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4010_ _4084_/B _4148_/C _4148_/D _4010_/D vssd2 vssd2 vccd2 vccd2 _4086_/B sky130_fd_sc_hd__or4_1
XFILLER_0_74_35 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5961_ _5962_/A _5962_/B _5962_/C vssd2 vssd2 vccd2 vccd2 _6059_/A sky130_fd_sc_hd__a21o_1
X_4912_ _4912_/A _4912_/B vssd2 vssd2 vccd2 vccd2 _4915_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__4634__D _4782_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_47_305 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7700_ _7798_/CLK _7700_/D vssd2 vssd2 vccd2 vccd2 _7700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_41 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5892_ _6550_/A _6812_/A vssd2 vssd2 vccd2 vccd2 _5915_/A sky130_fd_sc_hd__or2_1
X_7631_ _7641_/A vssd2 vssd2 vccd2 vccd2 _7631_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_114_85 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4843_ _4767_/A _4686_/A _4767_/B vssd2 vssd2 vccd2 vccd2 _4843_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_23_61 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6204__A _6707_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4774_ _4718_/A _4718_/B _4716_/X vssd2 vssd2 vccd2 vccd2 _4793_/A sky130_fd_sc_hd__o21ai_4
X_7562_ _7565_/A vssd2 vssd2 vccd2 vccd2 _7562_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_457 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_7_446 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6513_ _6590_/A _7294_/C vssd2 vssd2 vccd2 vccd2 _6515_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_55_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_43_544 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7493_ _7524_/A vssd2 vssd2 vccd2 vccd2 _7493_/Y sky130_fd_sc_hd__inv_2
X_6444_ _6445_/A _6445_/B vssd2 vssd2 vccd2 vccd2 _6444_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_70_396 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6375_ _6376_/A _6376_/B vssd2 vssd2 vccd2 vccd2 _6375_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_61_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4659__A _5468_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_11_441 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_23_290 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5326_ _5326_/A _5326_/B vssd2 vssd2 vccd2 vccd2 _5458_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_11_496 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5257_ _5257_/A _5257_/B vssd2 vssd2 vccd2 vccd2 _7747_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__6851__A1 _5991_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4208_ _4810_/A _4966_/A vssd2 vssd2 vccd2 vccd2 _4221_/A sky130_fd_sc_hd__nor2_1
X_5188_ _5119_/A _5119_/B _5117_/Y vssd2 vssd2 vccd2 vccd2 _5191_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_97_205 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4139_ _4139_/A _4193_/B vssd2 vssd2 vccd2 vccd2 _7730_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_249 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_78_430 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_65_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_38_338 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7829_ _7838_/CLK _7829_/D _7588_/Y vssd2 vssd2 vccd2 vccd2 _7829_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_444 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_19_552 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_93_488 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_34_522 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_34_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5342__B2 _5431_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout170 _6138_/A vssd2 vssd2 vccd2 vccd2 _6707_/A sky130_fd_sc_hd__clkbuf_8
Xfanout192 _4386_/X vssd2 vssd2 vccd2 vccd2 _4965_/B sky130_fd_sc_hd__clkbuf_8
Xfanout181 _6572_/B vssd2 vssd2 vccd2 vccd2 _7037_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_69_441 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_84_411 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_84_400 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1150 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_327 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1183 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_488 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__6024__A _6550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1194 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_56_157 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_71_127 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_37_382 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_37_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_107_281 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_52_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold618 _7812_/Q vssd2 vssd2 vccd2 vccd2 hold618/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold607 hold94/X vssd2 vssd2 vccd2 vccd2 _7873_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4490_ _4490_/A _4814_/B vssd2 vssd2 vccd2 vccd2 _4490_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_110_413 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_100_65 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold629 hold629/A vssd2 vssd2 vccd2 vccd2 hold629/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_569 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_901 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_260 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6160_ _6152_/X _6153_/X _6159_/X _5944_/B vssd2 vssd2 vccd2 vccd2 _7094_/A sky130_fd_sc_hd__o31a_4
XANTENNA__4629__D _5076_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_934 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _5111_/A _5111_/B vssd2 vssd2 vccd2 vccd2 _5114_/A sky130_fd_sc_hd__xor2_4
XTAP_923 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_282 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6091_ _6091_/A _6091_/B vssd2 vssd2 vccd2 vccd2 _6111_/A sky130_fd_sc_hd__xnor2_1
XTAP_978 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5097__B1 _5528_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_989 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _5042_/A _5042_/B _5374_/B _5528_/B vssd2 vssd2 vccd2 vccd2 _5043_/B sky130_fd_sc_hd__or4_1
XANTENNA__4926__B _4997_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6993_ _6357_/X _6359_/X _6281_/B _7143_/A vssd2 vssd2 vccd2 vccd2 _6995_/B sky130_fd_sc_hd__o211a_1
XANTENNA__4942__A _5207_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5944_ _6282_/A _5944_/B _5944_/C _5944_/D vssd2 vssd2 vccd2 vccd2 _5944_/X sky130_fd_sc_hd__and4_1
XFILLER_0_87_293 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5875_ _7844_/Q _6398_/B vssd2 vssd2 vccd2 vccd2 _5875_/X sky130_fd_sc_hd__and2_1
X_4826_ _4826_/A _4826_/B vssd2 vssd2 vccd2 vccd2 _4829_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_63_617 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA_fanout232_A _6588_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_16_500 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7614_ _7641_/A vssd2 vssd2 vccd2 vccd2 _7614_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_360 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_90_425 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_62_149 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7545_ _7561_/A vssd2 vssd2 vccd2 vccd2 _7545_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4757_ _4757_/A _4757_/B vssd2 vssd2 vccd2 vccd2 _4760_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_92 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6588__B _6588_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_43_385 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_43_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7476_ _7716_/Q _7483_/A2 _7483_/B1 hold337/X vssd2 vssd2 vccd2 vccd2 _7476_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_31_514 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4688_ _4618_/A _4619_/A _4618_/B vssd2 vssd2 vccd2 vccd2 _4688_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_113_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6427_ _6738_/A _6571_/C _6427_/C vssd2 vssd2 vccd2 vccd2 _6500_/B sky130_fd_sc_hd__and3_1
XFILLER_0_70_193 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4389__A _4962_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_3_460 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6358_ _6358_/A _6358_/B vssd2 vssd2 vccd2 vccd2 _6358_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_101_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5309_ _5257_/A _5256_/B _5548_/A vssd2 vssd2 vccd2 vccd2 _5310_/B sky130_fd_sc_hd__a21o_1
XANTENNA__6100__C _6282_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6289_ _6289_/A _6289_/B vssd2 vssd2 vccd2 vccd2 _6290_/B sky130_fd_sc_hd__xnor2_2
XPHY_200 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_21_wb_clk_i clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7776_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_222 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_211 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_81_469 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_34_330 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_34_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_34_385 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_104_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_34_396 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7403__A _7440_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4746__B _5528_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold4 hold4/A vssd2 vssd2 vccd2 vccd2 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6291__A2 _7047_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6043__A2 _5994_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_76_208 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6579__B1 _7099_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3990_ _3986_/X _3987_/X _3988_/X _3989_/X vssd2 vssd2 vccd2 vccd2 _3990_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_71_69 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_57_433 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_29_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_29_146 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_57_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_44_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5660_ _6019_/D _5979_/D vssd2 vssd2 vccd2 vccd2 _5662_/C sky130_fd_sc_hd__and2_1
X_4611_ _4539_/A _4539_/B _4537_/Y vssd2 vssd2 vccd2 vccd2 _4613_/B sky130_fd_sc_hd__a21boi_2
X_5591_ _5598_/B _5592_/C _7868_/Q vssd2 vssd2 vccd2 vccd2 _5594_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_44_149 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__5554__A1 _5528_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7330_ _7316_/A _7316_/B _7329_/X vssd2 vssd2 vccd2 vccd2 _7334_/D sky130_fd_sc_hd__a21oi_1
X_4542_ _4542_/A _4542_/B vssd2 vssd2 vccd2 vccd2 _4543_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6503__B1 _6430_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7261_ _7225_/A _7225_/B _7223_/B vssd2 vssd2 vccd2 vccd2 _7264_/B sky130_fd_sc_hd__a21oi_1
Xhold426 input32/X vssd2 vssd2 vccd2 vccd2 hold30/A sky130_fd_sc_hd__dlygate4sd3_1
X_4473_ _4474_/B _4474_/A vssd2 vssd2 vccd2 vccd2 _4473_/Y sky130_fd_sc_hd__nand2b_1
Xhold415 _7871_/Q vssd2 vssd2 vccd2 vccd2 hold415/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold404 _4049_/X vssd2 vssd2 vccd2 vccd2 hold404/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_536 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_13_558 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_110_221 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6212_ _6212_/A _6212_/B vssd2 vssd2 vccd2 vccd2 _6238_/A sky130_fd_sc_hd__xnor2_2
Xhold437 hold31/X vssd2 vssd2 vccd2 vccd2 input38/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 la_data_in[36] vssd2 vssd2 vccd2 vccd2 hold19/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 hold16/X vssd2 vssd2 vccd2 vccd2 _7841_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_265 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_96_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7192_ _7236_/A _7192_/B vssd2 vssd2 vccd2 vccd2 _7199_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__3868__A1 _7766_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6143_ _6144_/A _6144_/B vssd2 vssd2 vccd2 vccd2 _6199_/B sky130_fd_sc_hd__and2_1
XANTENNA__4937__A _5042_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_0_474 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_731 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _6074_/A _6253_/B _6253_/C _6191_/D vssd2 vssd2 vccd2 vccd2 _6078_/A sky130_fd_sc_hd__and4_1
X_5025_ _5072_/A _5025_/B vssd2 vssd2 vccd2 vccd2 _5027_/B sky130_fd_sc_hd__or2_2
XTAP_797 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA_fanout182_A _6103_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_45_70 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_67_219 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6590__C _7313_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6976_ _7037_/A _7291_/A _6977_/A vssd2 vssd2 vccd2 vccd2 _7040_/B sky130_fd_sc_hd__or3_1
XFILLER_0_48_400 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4045__A1 _4747_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4045__B2 _4598_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5927_ _6158_/A _6194_/C _6130_/C _6017_/B _7846_/Q vssd2 vssd2 vccd2 vccd2 _5927_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_63_403 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_48_488 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_48_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_90_233 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_75_285 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5858_ _5850_/B _5851_/X _5853_/X _5849_/X vssd2 vssd2 vccd2 vccd2 _5858_/X sky130_fd_sc_hd__a211o_1
X_5789_ _6071_/B _6019_/C _6019_/D vssd2 vssd2 vccd2 vccd2 _5826_/B sky130_fd_sc_hd__and3_1
X_4809_ _4809_/A _4809_/B vssd2 vssd2 vccd2 vccd2 _5164_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_90_277 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7528_ _7561_/A vssd2 vssd2 vccd2 vccd2 _7528_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_31_311 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7459_ _7699_/Q _7454_/C _7485_/B1 hold241/X vssd2 vssd2 vccd2 vccd2 _7459_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_31_344 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_31_366 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4847__A _5455_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_98_333 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_86_506 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6781__B _6939_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7369__S _7383_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_528 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_39_411 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5784__A1 _7844_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_39_433 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_81_222 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_81_211 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_499 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_54_458 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4339__A2 _4966_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5536__A1 _5468_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_10_528 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_66_58 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_89_366 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_106_53 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_82_68 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6830_ _6830_/A _6830_/B vssd2 vssd2 vccd2 vccd2 _6833_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_40 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_97 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6761_ _6763_/A _6763_/B vssd2 vssd2 vccd2 vccd2 _6762_/B sky130_fd_sc_hd__nand2_1
XANTENNA__6972__B1 _7313_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5712_ _5769_/B _6102_/B _6152_/C vssd2 vssd2 vccd2 vccd2 _5712_/X sky130_fd_sc_hd__and3b_1
X_3973_ _4125_/B _4022_/B vssd2 vssd2 vccd2 vccd2 _4057_/C sky130_fd_sc_hd__nor2_1
X_6692_ _6692_/A _6692_/B vssd2 vssd2 vccd2 vccd2 _6693_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_85_583 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5643_ _7856_/Q _7855_/Q _5645_/B vssd2 vssd2 vccd2 vccd2 _5644_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__5527__B2 _4814_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5574_ _5549_/A _5548_/B _5573_/X _5548_/A vssd2 vssd2 vccd2 vccd2 _7758_/D sky130_fd_sc_hd__a31oi_2
XFILLER_0_31_72 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7313_ _7313_/A _7313_/B vssd2 vssd2 vccd2 vccd2 _7313_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_53_491 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4525_ _5315_/B vssd2 vssd2 vccd2 vccd2 _4800_/C sky130_fd_sc_hd__inv_2
Xhold201 _7396_/X vssd2 vssd2 vccd2 vccd2 _7397_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_642 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold212 input88/X vssd2 vssd2 vccd2 vccd2 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _7467_/X vssd2 vssd2 vccd2 vccd2 _7707_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 hold373/X vssd2 vssd2 vccd2 vccd2 _7804_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_40_163 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_111_541 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold278 hold278/A vssd2 vssd2 vccd2 vccd2 la_data_out[10] sky130_fd_sc_hd__buf_12
Xhold267 hold620/X vssd2 vssd2 vccd2 vccd2 hold621/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 hold256/A vssd2 vssd2 vccd2 vccd2 la_data_out[0] sky130_fd_sc_hd__buf_12
X_7244_ _7244_/A _7244_/B vssd2 vssd2 vccd2 vccd2 _7246_/C sky130_fd_sc_hd__xnor2_1
Xhold245 _7738_/Q vssd2 vssd2 vccd2 vccd2 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ _4454_/Y _4455_/X _4103_/B vssd2 vssd2 vccd2 vccd2 _4456_/X sky130_fd_sc_hd__a21o_1
Xhold289 hold640/X vssd2 vssd2 vccd2 vccd2 hold641/A sky130_fd_sc_hd__dlygate4sd3_1
X_7175_ _7222_/A _7222_/B _7222_/C _7099_/B vssd2 vssd2 vccd2 vccd2 _7177_/A sky130_fd_sc_hd__a22o_1
XANTENNA__4667__A _4896_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4387_ _4810_/A _4965_/B vssd2 vssd2 vccd2 vccd2 _4391_/A sky130_fd_sc_hd__nor2_1
X_6126_ _6186_/A _6126_/B vssd2 vssd2 vccd2 vccd2 _6189_/B sky130_fd_sc_hd__nor2_1
XTAP_550 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ _6057_/A _6057_/B _6057_/C vssd2 vssd2 vccd2 vccd2 _6128_/A sky130_fd_sc_hd__and3_1
X_5008_ _5207_/A _5142_/C _5076_/D _5168_/A vssd2 vssd2 vccd2 vccd2 _5008_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5498__A _5498_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_76_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6959_ _6959_/A _6959_/B vssd2 vssd2 vccd2 vccd2 _6960_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_76_583 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_106_357 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6479__D _7051_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_182 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_32_675 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_563 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4577__A _5029_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_98_141 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_59_528 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4009__A1 _4809_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_52_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4009__B2 _4162_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_67_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_82_553 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_15_609 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_82_586 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_54_299 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_23_620 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_22_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5290_ _5217_/A _5217_/B _5215_/Y vssd2 vssd2 vccd2 vccd2 _5292_/B sky130_fd_sc_hd__a21bo_1
X_4310_ _4898_/A _4711_/A vssd2 vssd2 vccd2 vccd2 _4319_/B sky130_fd_sc_hd__or2_1
XFILLER_0_22_185 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_77_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4241_ _4242_/A _4243_/B vssd2 vssd2 vccd2 vccd2 _4303_/B sky130_fd_sc_hd__nor2_1
X_4172_ _5030_/A _5030_/B vssd2 vssd2 vccd2 vccd2 _4172_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4934__B _5404_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7862_ _7870_/CLK _7862_/D _7621_/Y vssd2 vssd2 vccd2 vccd2 _7862_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_58_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_58_550 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6813_ _6873_/A _7291_/A vssd2 vssd2 vccd2 vccd2 _6815_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_9_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5748__B2 _7844_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5748__A1 _7843_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7793_ _7793_/CLK _7793_/D _7552_/Y vssd2 vssd2 vccd2 vccd2 _7793_/Q sky130_fd_sc_hd__dfrtp_4
X_6744_ _6745_/B _6745_/A vssd2 vssd2 vccd2 vccd2 _6744_/X sky130_fd_sc_hd__and2b_1
X_3956_ _5030_/A vssd2 vssd2 vccd2 vccd2 _4729_/A sky130_fd_sc_hd__inv_2
XFILLER_0_85_391 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6675_ _6676_/A _6676_/B vssd2 vssd2 vccd2 vccd2 _6675_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_91_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_73_575 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_60_214 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5626_ _5581_/A _5581_/B _5645_/B vssd2 vssd2 vccd2 vccd2 _5632_/B sky130_fd_sc_hd__o21a_1
X_3887_ _4326_/C _4267_/D _4148_/B vssd2 vssd2 vccd2 vccd2 _3899_/D sky130_fd_sc_hd__nor3_1
XFILLER_0_33_417 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_103_305 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_103_349 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5557_ _5558_/A _5558_/B vssd2 vssd2 vccd2 vccd2 _5570_/A sky130_fd_sc_hd__nor2_1
X_4508_ _4810_/A _5222_/A _4462_/X _4464_/B vssd2 vssd2 vccd2 vccd2 _4516_/A sky130_fd_sc_hd__o31a_1
X_5488_ _5488_/A _5488_/B _5518_/B vssd2 vssd2 vccd2 vccd2 _5490_/A sky130_fd_sc_hd__and3_1
XANTENNA__6476__A2 _7222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7227_ _7259_/A _7227_/B vssd2 vssd2 vccd2 vccd2 _7229_/B sky130_fd_sc_hd__nand2_1
X_4439_ _4440_/A _4440_/B vssd2 vssd2 vccd2 vccd2 _4439_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_111_393 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5931__D _6664_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7158_ _7158_/A _7158_/B vssd2 vssd2 vccd2 vccd2 _7164_/A sky130_fd_sc_hd__xnor2_1
X_6109_ _6109_/A _6109_/B _6109_/C vssd2 vssd2 vccd2 vccd2 _6111_/B sky130_fd_sc_hd__nand3_1
X_7089_ _7153_/A _7089_/B vssd2 vssd2 vccd2 vccd2 _7109_/A sky130_fd_sc_hd__and2_1
XTAP_391 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5987__A1 _6157_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5987__B2 _7846_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1513 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XPHY_20 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_31 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XPHY_42 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_53 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_64 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_86 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_36_211 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_75 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_106_121 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_91_372 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_36_288 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_165 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_439 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_36_299 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5911__A1 _6402_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6787__A _7047_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4175__B1 _5029_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_20_656 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4100__A _4656_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6219__A2 _5816_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7411__A _7452_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_63_37 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6027__A _6138_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4790_ _4791_/A _4791_/B vssd2 vssd2 vccd2 vccd2 _4854_/A sky130_fd_sc_hd__and2_1
XFILLER_0_27_200 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3810_ _3831_/B _3811_/C _7802_/Q vssd2 vssd2 vccd2 vccd2 _3813_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_12_63 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_277 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6460_ _6313_/B _6313_/C _6385_/Y _6313_/A vssd2 vssd2 vccd2 vccd2 _6461_/B sky130_fd_sc_hd__a211o_1
X_6391_ _6390_/A _6390_/B _6390_/C vssd2 vssd2 vccd2 vccd2 _6392_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_556 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5411_ _5476_/A _5411_/B vssd2 vssd2 vccd2 vccd2 _5424_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_113_669 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xoutput125 hold661/X vssd2 vssd2 vccd2 vccd2 hold308/A sky130_fd_sc_hd__buf_6
Xoutput114 hold625/X vssd2 vssd2 vccd2 vccd2 hold274/A sky130_fd_sc_hd__buf_6
Xoutput103 hold667/X vssd2 vssd2 vccd2 vccd2 hold314/A sky130_fd_sc_hd__buf_6
X_5342_ _5394_/A _5341_/X _5207_/A _5431_/B vssd2 vssd2 vccd2 vccd2 _5344_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_11_612 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xoutput136 _7706_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[11] sky130_fd_sc_hd__buf_12
Xoutput158 _7726_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[31] sky130_fd_sc_hd__buf_12
Xoutput147 _7716_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[21] sky130_fd_sc_hd__buf_12
X_7012_ _7012_/A _7012_/B _7012_/C vssd2 vssd2 vccd2 vccd2 _7014_/A sky130_fd_sc_hd__or3_1
X_5273_ _5334_/B _5273_/B vssd2 vssd2 vccd2 vccd2 _5275_/B sky130_fd_sc_hd__nand2_1
X_4224_ _4088_/A _4088_/B _5029_/A vssd2 vssd2 vccd2 vccd2 _4226_/A sky130_fd_sc_hd__a21o_1
X_4155_ _4155_/A _4155_/B _4155_/C vssd2 vssd2 vccd2 vccd2 _5011_/A sky130_fd_sc_hd__and3_4
XFILLER_0_37_93 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4086_ _4814_/A _4086_/B vssd2 vssd2 vccd2 vccd2 _4087_/D sky130_fd_sc_hd__or2_1
XANTENNA__6630__A2 _7197_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7845_ _7854_/CLK _7845_/D _7604_/Y vssd2 vssd2 vccd2 vccd2 _7845_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6918__B1 _6669_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_65_328 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_108_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4988_ _4989_/A _4989_/B vssd2 vssd2 vccd2 vccd2 _4988_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_46_520 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7776_ _7776_/CLK _7776_/D _7535_/Y vssd2 vssd2 vccd2 vccd2 _7776_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_80_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4944__A2 _5276_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6727_ _6571_/B _7197_/A _6430_/B _6571_/A vssd2 vssd2 vccd2 vccd2 _6729_/A sky130_fd_sc_hd__a22o_1
X_3939_ _7779_/Q _7780_/Q _7781_/Q _3954_/C _4050_/B vssd2 vssd2 vccd2 vccd2 _3940_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_0_18_277 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6146__A1 _6664_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6146__B2 _5931_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6658_ _6658_/A _6658_/B vssd2 vssd2 vccd2 vccd2 _6660_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_383 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_61_523 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_18_299 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_103_113 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_14_450 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_258 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5609_ _5828_/B _5828_/C _5659_/B vssd2 vssd2 vccd2 vccd2 _6253_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_104_658 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6589_ _6590_/A _7313_/B vssd2 vssd2 vccd2 vccd2 _6591_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_61_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_14_472 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5016__A _5328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_88_409 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_68_122 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1332 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1354 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_177 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_56_306 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7377__S _7383_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1398 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_64_361 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_52_512 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_52_501 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__6137__A1 _5778_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xinput27 input27/A vssd2 vssd2 vccd2 vccd2 input27/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_236 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xinput16 input16/A vssd2 vssd2 vccd2 vccd2 input16/X sky130_fd_sc_hd__clkbuf_1
Xinput38 input38/A vssd2 vssd2 vccd2 vccd2 input38/X sky130_fd_sc_hd__clkbuf_1
Xinput49 wb_rst_i vssd2 vssd2 vccd2 vccd2 input49/X sky130_fd_sc_hd__buf_1
XFILLER_0_24_269 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_52_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_20_464 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_74_69 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5960_ _5960_/A _5960_/B vssd2 vssd2 vccd2 vccd2 _5962_/C sky130_fd_sc_hd__or2_1
XFILLER_0_59_100 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4911_ _4911_/A _4911_/B vssd2 vssd2 vccd2 vccd2 _4912_/B sky130_fd_sc_hd__xnor2_4
X_5891_ _6424_/A _6424_/B vssd2 vssd2 vccd2 vccd2 _6812_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_59_177 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7630_ _7641_/A vssd2 vssd2 vccd2 vccd2 _7630_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_114_53 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4842_ _4842_/A _4842_/B vssd2 vssd2 vccd2 vccd2 _4845_/A sky130_fd_sc_hd__and2_2
XANTENNA__5179__A2 _5550_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_23_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_114_97 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6204__B _6973_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4773_ _4920_/A _4773_/B vssd2 vssd2 vccd2 vccd2 _4834_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_62_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7561_ _7561_/A vssd2 vssd2 vccd2 vccd2 _7561_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_99_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4005__A _7765_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7492_ _7524_/A vssd2 vssd2 vccd2 vccd2 _7492_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_469 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6512_ _5744_/B _6510_/Y _6100_/D vssd2 vssd2 vccd2 vccd2 _7253_/C sky130_fd_sc_hd__a21o_4
X_6443_ _6369_/A _6369_/B _6367_/X vssd2 vssd2 vccd2 vccd2 _6445_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_15_247 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5887__B1 _6424_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6374_ _6299_/A _6299_/B _6297_/Y vssd2 vssd2 vccd2 vccd2 _6376_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_11_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5325_ _5325_/A _5498_/D vssd2 vssd2 vccd2 vccd2 _5330_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_54_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5256_ _5548_/A _5256_/B vssd2 vssd2 vccd2 vccd2 _5257_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5639__B1 _5645_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6851__A2 _5993_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4207_ _4199_/X _4200_/X _4206_/X _4080_/D vssd2 vssd2 vccd2 vccd2 _4207_/Y sky130_fd_sc_hd__o31ai_2
XANTENNA__4311__B1 _7771_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5187_ _5187_/A _5187_/B vssd2 vssd2 vccd2 vccd2 _5191_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__7051__A _7051_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4138_ _4189_/C _4138_/B vssd2 vssd2 vccd2 vccd2 _4193_/B sky130_fd_sc_hd__xnor2_1
X_4069_ _3986_/A _4125_/C _3986_/B _4067_/X _4068_/X vssd2 vssd2 vccd2 vccd2 _4069_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_65_103 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7828_ _7838_/CLK _7828_/D _7587_/Y vssd2 vssd2 vccd2 vccd2 _7828_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_456 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_65_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_46_350 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7759_ _7776_/CLK _7759_/D _7518_/Y vssd2 vssd2 vccd2 vccd2 _7759_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_34_512 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_28_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
Xfanout182 _6103_/X vssd2 vssd2 vccd2 vccd2 _7047_/A sky130_fd_sc_hd__buf_4
Xfanout193 _4386_/X vssd2 vssd2 vccd2 vccd2 _5328_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_57_604 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5802__B1 _6283_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1140 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_306 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XTAP_1173 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_136 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6024__B _6973_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1195 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4369__B1 _4782_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_44_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_37_361 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_71_139 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_64_180 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_52_320 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_4_417 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_107_293 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold608 _7807_/Q vssd2 vssd2 vccd2 vccd2 hold608/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_386 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold619 hold619/A vssd2 vssd2 vccd2 vccd2 hold619/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6975__A _7037_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6090_ _6090_/A _6090_/B vssd2 vssd2 vccd2 vccd2 _6091_/B sky130_fd_sc_hd__nand2_1
XTAP_935 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _5110_/A _5110_/B vssd2 vssd2 vccd2 vccd2 _5111_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_85_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_957 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5145_/A _5374_/B _5528_/B _5042_/A vssd2 vssd2 vccd2 vccd2 _5041_/X sky130_fd_sc_hd__o22a_1
XTAP_979 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_7 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_79_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
Xclkbuf_0_wb_clk_i wb_clk_i vssd2 vssd2 vccd2 vccd2 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_209 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6992_ _6281_/X _6284_/X _5937_/B _7143_/B vssd2 vssd2 vccd2 vccd2 _6995_/A sky130_fd_sc_hd__o211a_1
XFILLER_0_87_261 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4942__B _5366_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5943_ _5944_/B _5944_/C _5944_/D vssd2 vssd2 vccd2 vccd2 _5943_/X sky130_fd_sc_hd__and3_1
XANTENNA__6215__A _6812_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_47_136 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5874_ _6157_/A _6194_/C _6130_/C vssd2 vssd2 vccd2 vccd2 _5886_/A sky130_fd_sc_hd__and3_1
XFILLER_0_90_415 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_75_478 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4825_ _4825_/A _4825_/B vssd2 vssd2 vccd2 vccd2 _4826_/B sky130_fd_sc_hd__xnor2_4
X_7613_ _7613_/A vssd2 vssd2 vccd2 vccd2 _7613_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_62_106 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_47_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_90_437 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7544_ _7561_/A vssd2 vssd2 vccd2 vccd2 _7544_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_523 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_28_372 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_90_459 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4756_ _4756_/A _4756_/B vssd2 vssd2 vccd2 vccd2 _4757_/B sky130_fd_sc_hd__xor2_1
XANTENNA_fanout225_A _6549_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_180 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_16_556 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_71_673 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4687_ _4691_/A vssd2 vssd2 vccd2 vccd2 _4687_/Y sky130_fd_sc_hd__inv_2
X_7475_ _7715_/Q _7483_/A2 _7483_/B1 hold347/X vssd2 vssd2 vccd2 vccd2 _7475_/X sky130_fd_sc_hd__a22o_1
X_6426_ _6426_/A _6426_/B vssd2 vssd2 vccd2 vccd2 _6427_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__4389__B _5042_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_101_447 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6357_ _6510_/A _6357_/B vssd2 vssd2 vccd2 vccd2 _6357_/X sky130_fd_sc_hd__and2_2
X_5308_ _5308_/A _5308_/B vssd2 vssd2 vccd2 vccd2 _5357_/C sky130_fd_sc_hd__xnor2_4
X_6288_ _6590_/A _6289_/A _6430_/B vssd2 vssd2 vccd2 vccd2 _6288_/X sky130_fd_sc_hd__and3_1
X_5239_ _5239_/A _5239_/B vssd2 vssd2 vccd2 vccd2 _5240_/B sky130_fd_sc_hd__xnor2_4
XPHY_201 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_78_261 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_109_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XPHY_212 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_81_415 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_66_456 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_26_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_38_147 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_53_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_46_191 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_22_504 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_183 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4523__B1 _5458_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7390__S _7418_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold5 hold5/A vssd2 vssd2 vccd2 vccd2 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_526 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6579__A1 _6425_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6579__B2 _5931_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_72_404 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_29_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5003__A1 _5145_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_72_426 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4610_ _4610_/A _4610_/B vssd2 vssd2 vccd2 vccd2 _4613_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_489 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_44_117 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__5874__A _6157_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6736__D1 _7294_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_112_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_53_640 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5590_ _5645_/B _7867_/Q vssd2 vssd2 vccd2 vccd2 _5592_/C sky130_fd_sc_hd__and2_1
XFILLER_0_25_320 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5554__A2 _5431_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_37_191 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_4541_ _4542_/B _4542_/A vssd2 vssd2 vccd2 vccd2 _4541_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_80_492 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_481 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6503__A1 _6425_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7260_ _7289_/A _7260_/B vssd2 vssd2 vccd2 vccd2 _7267_/A sky130_fd_sc_hd__or2_1
X_4472_ _4350_/A _4350_/B _4408_/B _4409_/B _4409_/A vssd2 vssd2 vccd2 vccd2 _4474_/B
+ sky130_fd_sc_hd__a32oi_4
Xhold405 _7870_/Q vssd2 vssd2 vccd2 vccd2 _5821_/B sky130_fd_sc_hd__buf_2
Xhold427 hold30/X vssd2 vssd2 vccd2 vccd2 _7845_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 la_data_in[35] vssd2 vssd2 vccd2 vccd2 hold3/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_25_397 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6211_ _6212_/B _6212_/A vssd2 vssd2 vccd2 vccd2 _6261_/B sky130_fd_sc_hd__and2b_1
XANTENNA__6503__B2 _5931_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7191_ _7191_/A _7191_/B _7189_/Y vssd2 vssd2 vccd2 vccd2 _7192_/B sky130_fd_sc_hd__or3b_1
Xhold438 input38/X vssd2 vssd2 vccd2 vccd2 hold32/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 hold19/X vssd2 vssd2 vccd2 vccd2 input30/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_233 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6142_ _6142_/A _6142_/B vssd2 vssd2 vccd2 vccd2 _6144_/B sky130_fd_sc_hd__xnor2_2
XTAP_710 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_277 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4937__B _5550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_732 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7313__B _7313_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_776 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _6019_/D _6071_/X _6072_/X vssd2 vssd2 vccd2 vccd2 _6073_/Y sky130_fd_sc_hd__a21oi_2
X_5024_ _5024_/A _5024_/B _5024_/C vssd2 vssd2 vccd2 vccd2 _5025_/B sky130_fd_sc_hd__nor3_1
XTAP_798 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout175_A _4747_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_45_82 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_17_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5768__B _6550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6975_ _7037_/A _7291_/A vssd2 vssd2 vccd2 vccd2 _6977_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4045__A2 _4898_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5926_ _7844_/Q _5588_/Y _6398_/B _7845_/Q vssd2 vssd2 vccd2 vccd2 _5926_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_75_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_63_415 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_92 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5857_ _5857_/A _5857_/B _5857_/C _5857_/D vssd2 vssd2 vccd2 vccd2 _5857_/X sky130_fd_sc_hd__or4_1
XFILLER_0_90_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5788_ _5778_/X _5786_/Y _5736_/X vssd2 vssd2 vccd2 vccd2 _6636_/A sky130_fd_sc_hd__a21o_2
X_4808_ _4808_/A _4808_/B vssd2 vssd2 vccd2 vccd2 _4811_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_8_586 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_331 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_28_191 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_90_289 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4739_ _4739_/A _4739_/B vssd2 vssd2 vccd2 vccd2 _4749_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_150 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7527_ _7563_/A vssd2 vssd2 vccd2 vccd2 _7527_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_114_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7458_ _7698_/Q _7454_/C _7485_/B1 hold237/X vssd2 vssd2 vccd2 vccd2 _7458_/X sky130_fd_sc_hd__a22o_1
X_6409_ _6409_/A _6409_/B vssd2 vssd2 vccd2 vccd2 _6410_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_31_378 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7389_ _7440_/A _7389_/B vssd2 vssd2 vccd2 vccd2 _7663_/D sky130_fd_sc_hd__and2_1
XANTENNA__7470__A2 _7483_/A2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_98_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4863__A _4863_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6781__C _7253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5375__A2_N _5550_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_66_242 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_27_607 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_39_456 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_66_275 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_26_117 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5536__A2 _5431_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_105_572 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_62_492 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_22_323 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7461__A2 _7454_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5869__A _7336_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_77_529 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_65 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6760_ _6763_/A _6763_/B vssd2 vssd2 vccd2 vccd2 _6762_/A sky130_fd_sc_hd__or2_1
XFILLER_0_15_52 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6972__A1 _6571_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6972__B2 _6571_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5711_ _7877_/Q _5711_/B vssd2 vssd2 vccd2 vccd2 _5992_/B sky130_fd_sc_hd__xnor2_4
X_3972_ _4068_/B _4252_/B _4252_/D _4707_/A vssd2 vssd2 vccd2 vccd2 _4020_/B sky130_fd_sc_hd__nor4_2
X_6691_ _6692_/A _6692_/B vssd2 vssd2 vccd2 vccd2 _6691_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_57_286 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_45_426 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5642_ _6424_/A _5878_/B vssd2 vssd2 vccd2 vccd2 _5836_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_53_470 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5573_ _5570_/A _5570_/C _5573_/C _5573_/D vssd2 vssd2 vccd2 vccd2 _5573_/X sky130_fd_sc_hd__and4bb_1
X_7312_ _7326_/D _7312_/B vssd2 vssd2 vccd2 vccd2 _7834_/D sky130_fd_sc_hd__xnor2_1
Xhold202 hold369/X vssd2 vssd2 vccd2 vccd2 _7781_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4524_ _4519_/X _4520_/X _4523_/X _4458_/D vssd2 vssd2 vccd2 vccd2 _5414_/A sky130_fd_sc_hd__o31ai_4
Xhold235 _7733_/Q vssd2 vssd2 vccd2 vccd2 hold235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 _7416_/X vssd2 vssd2 vccd2 vccd2 _7417_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _7447_/X vssd2 vssd2 vccd2 vccd2 _7448_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_153 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_41_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_111_553 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
Xhold257 hold610/X vssd2 vssd2 vccd2 vccd2 hold611/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 hold268/A vssd2 vssd2 vccd2 vccd2 la_data_out[3] sky130_fd_sc_hd__buf_12
X_7243_ _7244_/A _7244_/B vssd2 vssd2 vccd2 vccd2 _7275_/B sky130_fd_sc_hd__and2b_1
Xhold246 _7466_/X vssd2 vssd2 vccd2 vccd2 _7706_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4455_ _3813_/A _3813_/B _4454_/B _3886_/C _3893_/B vssd2 vssd2 vccd2 vccd2 _4455_/X
+ sky130_fd_sc_hd__a2111o_1
X_7174_ _7174_/A _7326_/C vssd2 vssd2 vccd2 vccd2 _7830_/D sky130_fd_sc_hd__xnor2_1
Xhold279 hold630/X vssd2 vssd2 vccd2 vccd2 hold631/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4667__B _5220_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4386_ _4380_/Y _4382_/X _4385_/X _4144_/D vssd2 vssd2 vccd2 vccd2 _4386_/X sky130_fd_sc_hd__a31o_1
X_6125_ _6311_/A _6311_/B vssd2 vssd2 vccd2 vccd2 _6126_/B sky130_fd_sc_hd__and2_1
XTAP_540 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout292_A _7629_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_573 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _6055_/B _6055_/C _6055_/A vssd2 vssd2 vccd2 vccd2 _6057_/C sky130_fd_sc_hd__a21o_1
XTAP_595 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _4947_/A _4947_/B _4945_/Y vssd2 vssd2 vccd2 vccd2 _5027_/A sky130_fd_sc_hd__a21bo_2
XANTENNA__5498__B _5550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_95_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_72_80 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_48_220 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_76_551 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6958_ _6959_/A _6959_/B vssd2 vssd2 vccd2 vccd2 _6960_/A sky130_fd_sc_hd__and2_1
XFILLER_0_48_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5909_ _5909_/A _5909_/B vssd2 vssd2 vccd2 vccd2 _5910_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_286 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6889_ _6818_/Y _6822_/A _6932_/A _6888_/X vssd2 vssd2 vccd2 vccd2 _6891_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_91_565 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6715__A1 _6855_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4726__B1 _4880_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_63_267 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_51_429 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_17_673 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_32_643 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_102_575 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4577__B _4965_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_36_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_99_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_98_153 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_98_197 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6403__B1 _7051_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_39_220 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_82_521 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_67_595 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_54_201 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7409__A _7452_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_27_437 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_39_297 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_82_565 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_50_451 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_23_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_77_47 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4240_ _4243_/A _4242_/A _4243_/B vssd2 vssd2 vccd2 vccd2 _4244_/A sky130_fd_sc_hd__and3_1
X_4171_ _4171_/A _4171_/B _4171_/C _4171_/D vssd2 vssd2 vccd2 vccd2 _5030_/B sky130_fd_sc_hd__or4_4
XFILLER_0_93_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5996__A2 _5948_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_26_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__5599__A _7842_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_26_62 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7861_ _7870_/CLK _7861_/D _7620_/Y vssd2 vssd2 vccd2 vccd2 _7861_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6207__B _7037_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6812_ _6812_/A _6812_/B _7253_/C _7253_/D vssd2 vssd2 vccd2 vccd2 _6815_/B sky130_fd_sc_hd__or4_1
XFILLER_0_92_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5748__A2 _6281_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7792_ _7793_/CLK _7792_/D _7551_/Y vssd2 vssd2 vccd2 vccd2 _7792_/Q sky130_fd_sc_hd__dfrtp_4
X_6743_ _6677_/A _6677_/B _6675_/Y vssd2 vssd2 vccd2 vccd2 _6745_/B sky130_fd_sc_hd__o21a_1
X_3955_ _3955_/A _3955_/B vssd2 vssd2 vccd2 vccd2 _5030_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_42_50 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_73_532 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6674_ _6668_/A _7222_/B _6592_/B _6590_/X vssd2 vssd2 vccd2 vccd2 _6676_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_42_72 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3886_ _4457_/B _4519_/C _3886_/C vssd2 vssd2 vccd2 vccd2 _3886_/X sky130_fd_sc_hd__and3_1
X_5625_ _6191_/D _5630_/B _6075_/C vssd2 vssd2 vccd2 vccd2 _5655_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_84_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_5_353 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_317 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5556_ _5556_/A _5556_/B vssd2 vssd2 vccd2 vccd2 _5558_/B sky130_fd_sc_hd__xnor2_1
X_4507_ _4449_/A _4449_/B _4447_/Y vssd2 vssd2 vccd2 vccd2 _4517_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__5781__B _5781_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5487_ _5487_/A _5487_/B vssd2 vssd2 vccd2 vccd2 _5518_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_361 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7226_ _7145_/A _7313_/B _6669_/X _7143_/B vssd2 vssd2 vccd2 vccd2 _7227_/B sky130_fd_sc_hd__a22o_1
X_4438_ _4438_/A _4438_/B vssd2 vssd2 vccd2 vccd2 _4440_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__4397__B _5030_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7157_ _7158_/A _7158_/B vssd2 vssd2 vccd2 vccd2 _7157_/X sky130_fd_sc_hd__or2_1
X_4369_ _4863_/A _4711_/A _4782_/B _4898_/A vssd2 vssd2 vccd2 vccd2 _4370_/C sky130_fd_sc_hd__o22a_1
X_6108_ _6045_/A _6045_/B _6045_/C vssd2 vssd2 vccd2 vccd2 _6109_/C sky130_fd_sc_hd__a21bo_1
X_7088_ _6657_/B _7313_/B _6669_/X _6571_/B vssd2 vssd2 vccd2 vccd2 _7089_/B sky130_fd_sc_hd__a22o_1
XTAP_392 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6633__B1 _7253_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6039_ _6510_/A _5769_/X _5943_/X _6093_/A _6038_/X vssd2 vssd2 vccd2 vccd2 _6039_/X
+ sky130_fd_sc_hd__a221o_4
XANTENNA__5987__A2 _6281_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1503 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_90 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_68_348 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_21 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_10 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XPHY_32 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_43 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_54 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_65 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1569 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_87 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_76 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_64_587 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_106_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_51_237 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_177 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6787__B _7094_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6872__B1 _7313_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_99_462 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_87_602 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5212__A _5276_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6027__B _6812_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_101 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_59_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_86_178 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_55_532 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_12_97 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_113_626 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_113_615 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6390_ _6390_/A _6390_/B _6390_/C vssd2 vssd2 vccd2 vccd2 _6392_/A sky130_fd_sc_hd__and3_1
XFILLER_0_70_568 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5410_ _5475_/A _5475_/B vssd2 vssd2 vccd2 vccd2 _5411_/B sky130_fd_sc_hd__nand2_1
Xoutput115 hold655/X vssd2 vssd2 vccd2 vccd2 hold302/A sky130_fd_sc_hd__buf_6
Xoutput104 hold649/X vssd2 vssd2 vccd2 vccd2 hold296/A sky130_fd_sc_hd__buf_6
X_5341_ _5341_/A _5341_/B _5341_/C vssd2 vssd2 vccd2 vccd2 _5341_/X sky130_fd_sc_hd__or3_1
XFILLER_0_100_309 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xoutput126 hold621/X vssd2 vssd2 vccd2 vccd2 hold268/A sky130_fd_sc_hd__buf_6
Xoutput137 _7707_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[12] sky130_fd_sc_hd__buf_12
Xoutput159 _7698_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[3] sky130_fd_sc_hd__buf_12
Xoutput148 _7717_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[22] sky130_fd_sc_hd__buf_12
X_7011_ _7077_/A _7010_/X _6939_/A _7291_/B vssd2 vssd2 vccd2 vccd2 _7012_/C sky130_fd_sc_hd__o2bb2a_1
X_5272_ _5272_/A _5272_/B vssd2 vssd2 vccd2 vccd2 _5273_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5666__A1 _6282_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4223_ _4729_/A _4898_/A _5030_/B vssd2 vssd2 vccd2 vccd2 _4228_/A sky130_fd_sc_hd__or3b_1
XANTENNA__7602__A _7627_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4154_ _4081_/C _4101_/Y _4153_/X _4004_/B vssd2 vssd2 vccd2 vccd2 _4155_/C sky130_fd_sc_hd__a22oi_2
XANTENNA__6218__A _6668_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4085_ _4002_/Y _4084_/X _4083_/X vssd2 vssd2 vccd2 vccd2 _4087_/C sky130_fd_sc_hd__o21ba_1
XFILLER_0_78_602 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_77_134 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA_fanout255_A _6253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7844_ _7854_/CLK _7844_/D _7603_/Y vssd2 vssd2 vccd2 vccd2 _7844_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6918__B2 _6664_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6918__A1 _6738_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_77_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_53_93 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7775_ _7779_/CLK _7775_/D _7534_/Y vssd2 vssd2 vccd2 vccd2 _7775_/Q sky130_fd_sc_hd__dfrtp_4
X_4987_ _4916_/A _4916_/B _4914_/Y vssd2 vssd2 vccd2 vccd2 _4989_/B sky130_fd_sc_hd__a21oi_4
X_6726_ _6667_/A _6667_/B _6664_/X vssd2 vssd2 vccd2 vccd2 _6733_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_46_554 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3938_ _7779_/Q _7780_/Q _3954_/C _4050_/B vssd2 vssd2 vccd2 vccd2 _3944_/B sky130_fd_sc_hd__o31a_2
XANTENNA__6146__A2 _5948_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6657_ _7047_/A _6657_/B vssd2 vssd2 vccd2 vccd2 _6658_/B sky130_fd_sc_hd__and2_1
XFILLER_0_61_535 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3869_ _4457_/B _4519_/C _3868_/X _4656_/C _7760_/Q vssd2 vssd2 vccd2 vccd2 _3869_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5792__A _7845_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_33_204 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_104_637 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6588_ _6670_/A _6588_/B vssd2 vssd2 vccd2 vccd2 _7253_/D sky130_fd_sc_hd__nand2_2
X_5608_ _5828_/B _5828_/C vssd2 vssd2 vccd2 vccd2 _5608_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_103_125 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_14_484 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5539_ _5539_/A _5539_/B _5539_/C vssd2 vssd2 vccd2 vccd2 _5540_/B sky130_fd_sc_hd__or3_1
XFILLER_0_103_169 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4201__A _4809_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7209_ _7209_/A _7209_/B vssd2 vssd2 vccd2 vccd2 _7210_/B sky130_fd_sc_hd__or2_1
XANTENNA__5016__B _5366_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_wb_clk_i clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7802_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__7512__A _7564_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_96_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1322 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_159 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_91_181 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6137__A2 _5786_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xinput17 input17/A vssd2 vssd2 vccd2 vccd2 input17/X sky130_fd_sc_hd__clkbuf_1
Xinput28 input28/A vssd2 vssd2 vccd2 vccd2 input28/X sky130_fd_sc_hd__clkbuf_1
Xinput39 input39/A vssd2 vssd2 vccd2 vccd2 input39/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_248 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5207__A _5207_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_20_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_20_443 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_20_454 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4320__A1 _4598_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7422__A _7440_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_74_59 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_99_281 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_87_443 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4910_ _4911_/A _4911_/B vssd2 vssd2 vccd2 vccd2 _4910_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_59_145 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5890_ _5890_/A _5890_/B vssd2 vssd2 vccd2 vccd2 _5931_/C sky130_fd_sc_hd__or2_4
XFILLER_0_87_465 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4841_ _4841_/A _4841_/B vssd2 vssd2 vccd2 vccd2 _4842_/B sky130_fd_sc_hd__or2_1
XFILLER_0_47_318 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_75_649 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4772_ _4772_/A _4772_/B _4770_/Y vssd2 vssd2 vccd2 vccd2 _4773_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_43_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_7_426 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7560_ _7561_/A vssd2 vssd2 vccd2 vccd2 _7560_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_513 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7491_ _7524_/A vssd2 vssd2 vccd2 vccd2 _7491_/Y sky130_fd_sc_hd__inv_2
X_6511_ _5744_/B _6510_/Y _6100_/D vssd2 vssd2 vccd2 vccd2 _7294_/C sky130_fd_sc_hd__a21oi_4
XFILLER_0_28_587 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6442_ _6442_/A _6442_/B vssd2 vssd2 vccd2 vccd2 _6445_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_568 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_70_376 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_70_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6373_ _6373_/A _6373_/B vssd2 vssd2 vccd2 vccd2 _6376_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5324_ _5324_/A _5324_/B vssd2 vssd2 vccd2 vccd2 _5336_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_465 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4021__A _4328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_11_487 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5255_ _5357_/A _5357_/B vssd2 vssd2 vccd2 vccd2 _5256_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_47_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4206_ _4206_/A _4206_/B _4206_/C _4206_/D vssd2 vssd2 vccd2 vccd2 _4206_/X sky130_fd_sc_hd__or4_1
X_5186_ _5186_/A _5186_/B vssd2 vssd2 vccd2 vccd2 _5187_/B sky130_fd_sc_hd__xor2_2
XANTENNA__7051__B _7224_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4137_ _4189_/A _4187_/A vssd2 vssd2 vccd2 vccd2 _4138_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_78_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4068_ _7762_/Q _4068_/B vssd2 vssd2 vccd2 vccd2 _4068_/X sky130_fd_sc_hd__and2_1
X_7827_ _7838_/CLK _7827_/D _7586_/Y vssd2 vssd2 vccd2 vccd2 _7827_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_498 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_78_465 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_19_532 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_93_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7758_ _7758_/CLK _7758_/D _7517_/Y vssd2 vssd2 vccd2 vccd2 _7758_/Q sky130_fd_sc_hd__dfrtp_1
X_6709_ _6039_/X _6040_/X _7143_/B _5992_/B vssd2 vssd2 vccd2 vccd2 _6712_/A sky130_fd_sc_hd__o211a_1
XFILLER_0_46_384 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7689_ _7802_/CLK _7689_/D vssd2 vssd2 vccd2 vccd2 _7689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_434 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4866__A _5210_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout183 _6103_/X vssd2 vssd2 vccd2 vccd2 _6571_/C sky130_fd_sc_hd__clkbuf_2
Xfanout172 _6150_/A vssd2 vssd2 vccd2 vccd2 _6668_/A sky130_fd_sc_hd__buf_4
Xfanout194 _5325_/A vssd2 vssd2 vccd2 vccd2 _5220_/A sky130_fd_sc_hd__buf_4
XANTENNA__5263__C1 _4267_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7388__S _7418_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_96_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1141 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1196 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4369__B2 _4898_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4369__A1 _4863_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_25_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_25_513 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_25_535 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_114_209 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_107_261 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_64_192 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_4_429 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7417__A _7450_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_80_674 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xhold609 hold609/A vssd2 vssd2 vccd2 vccd2 hold609/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_527 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6975__B _7291_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_925 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5220_/A _5222_/A vssd2 vssd2 vccd2 vccd2 _5044_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_85_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_969 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_18_52 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_79_229 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6991_ _6991_/A _6991_/B vssd2 vssd2 vccd2 vccd2 _7001_/A sky130_fd_sc_hd__xnor2_1
X_5942_ _6093_/A _5992_/B _5992_/C vssd2 vssd2 vccd2 vccd2 _5947_/C sky130_fd_sc_hd__and3_1
XFILLER_0_87_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_34_73 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6215__B _6812_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_75_446 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_75_435 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5873_ _7845_/Q _6017_/B vssd2 vssd2 vccd2 vccd2 _5873_/X sky130_fd_sc_hd__and2_1
XFILLER_0_90_405 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4824_ _4825_/A _4825_/B vssd2 vssd2 vccd2 vccd2 _4824_/Y sky130_fd_sc_hd__nand2b_1
X_7612_ _7613_/A vssd2 vssd2 vccd2 vccd2 _7612_/Y sky130_fd_sc_hd__inv_2
X_4755_ _4756_/A _4756_/B vssd2 vssd2 vccd2 vccd2 _4755_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_62_118 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7543_ _7561_/A vssd2 vssd2 vccd2 vccd2 _7543_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_384 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5309__B1 _5548_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4686_ _4686_/A _4686_/B vssd2 vssd2 vccd2 vccd2 _4691_/A sky130_fd_sc_hd__and2_2
X_7474_ _7714_/Q _7483_/A2 _7483_/B1 hold333/X vssd2 vssd2 vccd2 vccd2 _7474_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_31_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA_fanout218_A _4628_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5129__A1_N _4996_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6425_ _6425_/A _7094_/A _6426_/B vssd2 vssd2 vccd2 vccd2 _6500_/A sky130_fd_sc_hd__and3_1
X_6356_ _5816_/A _5816_/B _7237_/A vssd2 vssd2 vccd2 vccd2 _6364_/A sky130_fd_sc_hd__a21oi_2
X_5307_ _5254_/A _5254_/B _5247_/A vssd2 vssd2 vccd2 vccd2 _5308_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_11_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6287_ _6590_/A _6430_/B vssd2 vssd2 vccd2 vccd2 _6289_/B sky130_fd_sc_hd__nand2_1
XANTENNA__7482__B1 _7483_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5238_ _5239_/B _5239_/A vssd2 vssd2 vccd2 vccd2 _5238_/X sky130_fd_sc_hd__and2b_1
X_5169_ _5169_/A _5169_/B vssd2 vssd2 vccd2 vccd2 _5171_/B sky130_fd_sc_hd__xor2_1
XANTENNA__5310__A _5357_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6993__C1 _7143_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_38_104 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_224 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_213 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_202 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_38_137 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_109_515 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_81_405 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_81_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_74_490 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7237__A _7237_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_104_253 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_22_538 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__7473__B1 _7483_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_100_481 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xhold6 hold6/A vssd2 vssd2 vccd2 vccd2 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6579__A2 _6430_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4039__B1 _7761_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5787__B1 _5736_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_240 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_57_402 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5220__A _5220_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_57_446 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6035__B _6281_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_57_457 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6736__C1 _7222_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_29_159 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5003__A2 _5404_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_72_438 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_72_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_111_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_105_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4540_ _4407_/A _4407_/B _4470_/B _4471_/B _4471_/A vssd2 vssd2 vccd2 vccd2 _4542_/B
+ sky130_fd_sc_hd__a32oi_4
XANTENNA__6503__A2 _7197_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold406 _5820_/X vssd2 vssd2 vccd2 vccd2 _6069_/A sky130_fd_sc_hd__buf_2
X_4471_ _4471_/A _4471_/B vssd2 vssd2 vccd2 vccd2 _4474_/A sky130_fd_sc_hd__xor2_2
Xhold417 hold3/X vssd2 vssd2 vccd2 vccd2 input29/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_387 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6210_ _6210_/A _6210_/B vssd2 vssd2 vccd2 vccd2 _6212_/B sky130_fd_sc_hd__xnor2_2
Xhold439 hold32/X vssd2 vssd2 vccd2 vccd2 _7850_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7190_ _7191_/A _7191_/B _7232_/B _7189_/B vssd2 vssd2 vccd2 vccd2 _7236_/A sky130_fd_sc_hd__o211a_1
Xhold428 la_data_in[10] vssd2 vssd2 vccd2 vccd2 hold5/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6141_ _6142_/B _6142_/A vssd2 vssd2 vccd2 vccd2 _6199_/A sky130_fd_sc_hd__and2b_1
XTAP_700 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_289 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_0_465 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_29_40 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_29_62 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_722 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7464__B1 _7485_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_29_84 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6072_ _6282_/A _6016_/B _6071_/B _6017_/B _7849_/Q vssd2 vssd2 vccd2 vccd2 _6072_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_744 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _5024_/A _5024_/B _5024_/C vssd2 vssd2 vccd2 vccd2 _5072_/A sky130_fd_sc_hd__o21a_1
XTAP_799 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7610__A _7613_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_45_61 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_45_50 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA_fanout168_A _6215_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6974_ _6974_/A _7040_/A vssd2 vssd2 vccd2 vccd2 _6977_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_210 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_48_413 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5925_ _7847_/Q _6016_/B _6071_/B vssd2 vssd2 vccd2 vccd2 _5925_/X sky130_fd_sc_hd__and3_1
X_5856_ _6283_/A _5936_/B _5936_/C vssd2 vssd2 vccd2 vccd2 _5857_/D sky130_fd_sc_hd__and3_1
X_4807_ _4807_/A _4880_/B vssd2 vssd2 vccd2 vccd2 _4808_/B sky130_fd_sc_hd__or2_2
XFILLER_0_61_71 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_507 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5787_ _5778_/X _5786_/Y _5736_/X vssd2 vssd2 vccd2 vccd2 _6082_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_63_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5950__B1 _5948_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4738_ _4739_/A _4739_/B vssd2 vssd2 vccd2 vccd2 _4738_/Y sky130_fd_sc_hd__nand2b_1
X_7526_ _7561_/A vssd2 vssd2 vccd2 vccd2 _7526_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_114_551 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4669_ _4669_/A _4669_/B vssd2 vssd2 vccd2 vccd2 _4670_/B sky130_fd_sc_hd__xnor2_1
X_7457_ _7697_/Q _7454_/C _7485_/B1 hold247/X vssd2 vssd2 vccd2 vccd2 _7457_/X sky130_fd_sc_hd__a22o_1
X_6408_ _6409_/A _6409_/B vssd2 vssd2 vccd2 vccd2 _6408_/X sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_101_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7388_ hold153/X _7775_/D _7418_/S vssd2 vssd2 vccd2 vccd2 _7388_/X sky130_fd_sc_hd__mux2_1
X_6339_ _6276_/A _6276_/B _6276_/C vssd2 vssd2 vccd2 vccd2 _6347_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__4269__B1 _7766_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7455__B1 _7485_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5006__A1_N _4863_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7520__A _7557_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4863__B _5550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6781__D _7253_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6136__A _6550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_519 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5040__A _5220_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_94_563 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_66_232 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_39_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_41_19 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_54_438 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_54_416 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_479 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_50_600 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_22_302 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_105_551 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_62_471 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_22_313 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7430__A _7436_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_89_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_82_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_82_59 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_106_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_3971_ _3971_/A vssd2 vssd2 vccd2 vccd2 _3971_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4432__B1 _4782_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_57_243 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6972__A2 _7294_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5710_ _7878_/Q _5710_/B vssd2 vssd2 vccd2 vccd2 _5769_/B sky130_fd_sc_hd__xor2_4
X_6690_ _6608_/A _6608_/B _6606_/Y vssd2 vssd2 vccd2 vccd2 _6692_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_72_213 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_72_202 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6709__C1 _5992_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_57_298 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_45_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5641_ _7859_/Q _5641_/B vssd2 vssd2 vccd2 vccd2 _5878_/B sky130_fd_sc_hd__xor2_4
XANTENNA__5932__B1 _6812_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_60_408 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5572_ _5572_/A _5572_/B vssd2 vssd2 vccd2 vccd2 _7756_/D sky130_fd_sc_hd__xnor2_1
X_7311_ _7219_/B _7335_/A _6069_/A vssd2 vssd2 vccd2 vccd2 _7312_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_13_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4523_ _4521_/Y _4522_/X _5458_/A vssd2 vssd2 vccd2 vccd2 _4523_/X sky130_fd_sc_hd__o21a_1
X_7242_ _7242_/A _7242_/B vssd2 vssd2 vccd2 vccd2 _7244_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__7605__A _7627_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold203 _7400_/X vssd2 vssd2 vccd2 vccd2 _7401_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 hold399/X vssd2 vssd2 vccd2 vccd2 _7794_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 hold356/X vssd2 vssd2 vccd2 vccd2 _7805_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 hold258/A vssd2 vssd2 vccd2 vccd2 la_data_out[7] sky130_fd_sc_hd__buf_12
Xhold269 hold622/X vssd2 vssd2 vccd2 vccd2 hold623/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _7729_/Q vssd2 vssd2 vccd2 vccd2 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 _7461_/X vssd2 vssd2 vccd2 vccd2 _7701_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ _4454_/A _4454_/B vssd2 vssd2 vccd2 vccd2 _4454_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_40_176 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7173_ _7211_/D _7173_/B vssd2 vssd2 vccd2 vccd2 _7326_/C sky130_fd_sc_hd__xor2_4
X_4385_ _4706_/A1 _4075_/B _4384_/Y _4809_/B vssd2 vssd2 vccd2 vccd2 _4385_/X sky130_fd_sc_hd__o2bb2a_1
X_6124_ _6311_/A _6311_/B vssd2 vssd2 vccd2 vccd2 _6186_/A sky130_fd_sc_hd__nor2_1
XTAP_530 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6055_/A _6055_/B _6055_/C vssd2 vssd2 vccd2 vccd2 _6057_/B sky130_fd_sc_hd__nand3_1
XTAP_574 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _4863_/A _5431_/B _5123_/A _5005_/Y vssd2 vssd2 vccd2 vccd2 _5060_/A sky130_fd_sc_hd__a2bb2o_2
XANTENNA_fanout285_A _7564_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_596 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_305 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5498__C _5528_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6957_ _6891_/A _6891_/C _6891_/B vssd2 vssd2 vccd2 vccd2 _6959_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__4423__B1 _5455_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5795__A _7846_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5908_ _5908_/A vssd2 vssd2 vccd2 vccd2 _5909_/B sky130_fd_sc_hd__inv_2
XFILLER_0_63_202 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6888_ _6887_/A _6887_/B _6875_/X vssd2 vssd2 vccd2 vccd2 _6888_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__4650__C_N _5030_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6715__A2 _7181_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5839_ _6093_/A _5878_/B _5878_/C vssd2 vssd2 vccd2 vccd2 _5839_/X sky130_fd_sc_hd__and3_1
XFILLER_0_8_351 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_8_340 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4204__A _7766_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_44_493 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7509_ _7565_/A vssd2 vssd2 vccd2 vccd2 _7509_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_102_510 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__7515__A _7564_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_31_187 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_587 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5151__A1 _5276_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_98_121 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_98_165 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6403__B2 _6707_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6403__A1 _6783_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_316 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_52_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_67_541 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7396__S _7418_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_82_511 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_27_405 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_39_265 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_27_449 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_82_577 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_54_257 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_112_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_77_15 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_50_463 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_4170_ _4706_/A1 _4029_/X _4030_/X _7767_/Q _4169_/X vssd2 vssd2 vccd2 vccd2 _4171_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4784__A _4966_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_93_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7860_ _7886_/CLK _7860_/D _7619_/Y vssd2 vssd2 vccd2 vccd2 _7860_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_74 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_77_327 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6811_ _5890_/A _5890_/B _6664_/A _7294_/C _7313_/B vssd2 vssd2 vccd2 vccd2 _6811_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_26_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7791_ _7795_/CLK _7791_/D _7550_/Y vssd2 vssd2 vccd2 vccd2 _7791_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6504__A _6812_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6742_ _6742_/A _6742_/B vssd2 vssd2 vccd2 vccd2 _6745_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_574 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3954_ _4050_/B _7779_/Q _3954_/C vssd2 vssd2 vccd2 vccd2 _3955_/B sky130_fd_sc_hd__and3_1
XFILLER_0_85_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_73_544 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6673_ _6673_/A _6673_/B vssd2 vssd2 vccd2 vccd2 _6676_/A sky130_fd_sc_hd__xor2_2
X_3885_ _3813_/A _3813_/B _4745_/A _4454_/B _3830_/X vssd2 vssd2 vccd2 vccd2 _4149_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_60_205 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4024__A _4893_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5624_ _6253_/B _6253_/C _5617_/X _7313_/A _7840_/Q vssd2 vssd2 vccd2 vccd2 _5624_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_26_460 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_103_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5555_ _5537_/A _5537_/B _5534_/X vssd2 vssd2 vccd2 vccd2 _5556_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__3863__A _4268_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_77_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4506_ _4506_/A _4506_/B vssd2 vssd2 vccd2 vccd2 _4539_/A sky130_fd_sc_hd__xnor2_2
X_5486_ _5486_/A _5486_/B _5487_/A vssd2 vssd2 vccd2 vccd2 _5486_/X sky130_fd_sc_hd__and3_1
X_7225_ _7225_/A _7225_/B vssd2 vssd2 vccd2 vccd2 _7229_/A sky130_fd_sc_hd__xnor2_1
X_4437_ _4438_/A _4438_/B vssd2 vssd2 vccd2 vccd2 _4506_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_111_373 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7156_ _7154_/Y _7155_/X _7037_/A _6670_/Y vssd2 vssd2 vccd2 vccd2 _7158_/B sky130_fd_sc_hd__o2bb2a_1
XANTENNA__4397__C _5030_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6107_ _6106_/B _6106_/C _6106_/A vssd2 vssd2 vccd2 vccd2 _6109_/B sky130_fd_sc_hd__a21o_1
X_4368_ _4367_/B _4438_/A vssd2 vssd2 vccd2 vccd2 _4441_/A sky130_fd_sc_hd__and2b_2
XTAP_360 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7087_ _7087_/A _7087_/B vssd2 vssd2 vccd2 vccd2 _7828_/D sky130_fd_sc_hd__xnor2_1
XTAP_393 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _4299_/A _4299_/B vssd2 vssd2 vccd2 vccd2 _4303_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__6633__B2 _6707_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6633__A1 _6783_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6038_ _7846_/Q _6510_/B _5992_/C _6253_/A vssd2 vssd2 vccd2 vccd2 _6038_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_68_305 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_22 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_11 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_552 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_49_541 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_33 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_44 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_308 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XPHY_88 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_66 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_76_382 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_99 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_36_224 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_91_341 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_36_268 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6787__C _7143_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_32_441 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_20_614 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6872__A1 _6424_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6872__B2 _6664_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_63_17 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5212__B _5406_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_99_474 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_87_669 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_55_511 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_12_43 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_27_257 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_268 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_70_525 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_15_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_42_216 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4779__A _4779_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xoutput116 hold659/X vssd2 vssd2 vccd2 vccd2 hold306/A sky130_fd_sc_hd__buf_6
Xoutput105 hold635/X vssd2 vssd2 vccd2 vccd2 hold282/A sky130_fd_sc_hd__buf_6
X_5340_ _5341_/A _5341_/B _5341_/C vssd2 vssd2 vccd2 vccd2 _5394_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_23_463 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xoutput127 hold617/X vssd2 vssd2 vccd2 vccd2 hold264/A sky130_fd_sc_hd__buf_6
X_5271_ _5272_/A _5272_/B vssd2 vssd2 vccd2 vccd2 _5334_/B sky130_fd_sc_hd__or2_1
Xoutput138 _7708_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[13] sky130_fd_sc_hd__buf_12
Xoutput149 _7718_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[23] sky130_fd_sc_hd__buf_12
XANTENNA__6863__A1 _6150_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7010_ _7010_/A _7010_/B _7008_/X vssd2 vssd2 vccd2 vccd2 _7010_/X sky130_fd_sc_hd__or3b_1
X_4222_ _4178_/A _4178_/B _4176_/Y vssd2 vssd2 vccd2 vccd2 _4232_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_179 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4153_ _4809_/A _4002_/A _4002_/B _4002_/C _4152_/X vssd2 vssd2 vccd2 vccd2 _4153_/X
+ sky130_fd_sc_hd__a41o_1
X_4084_ _4457_/A _4084_/B _4004_/B vssd2 vssd2 vccd2 vccd2 _4084_/X sky130_fd_sc_hd__or3b_1
XANTENNA__6218__B _7047_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_77_102 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_78_658 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7843_ _7854_/CLK _7843_/D _7602_/Y vssd2 vssd2 vccd2 vccd2 _7843_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6918__A2 _7313_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_93_617 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4986_ _4986_/A _4986_/B vssd2 vssd2 vccd2 vccd2 _4989_/A sky130_fd_sc_hd__xnor2_4
X_7774_ _7806_/CLK _7774_/D _7533_/Y vssd2 vssd2 vccd2 vccd2 _7774_/Q sky130_fd_sc_hd__dfrtp_1
X_6725_ _6656_/A _6658_/B _6656_/B vssd2 vssd2 vccd2 vccd2 _6734_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_46_544 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_46_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3937_ _4022_/B _4162_/B vssd2 vssd2 vccd2 vccd2 _4315_/C sky130_fd_sc_hd__nor2_1
XANTENNA_fanout248_A _4809_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_46_566 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_104_605 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6656_ _6656_/A _6656_/B vssd2 vssd2 vccd2 vccd2 _6658_/A sky130_fd_sc_hd__nand2_1
X_3868_ _7766_/Q _4326_/B _4326_/C _7764_/Q _4458_/D vssd2 vssd2 vccd2 vccd2 _3868_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_61_569 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6587_ _6587_/A _6587_/B vssd2 vssd2 vccd2 vccd2 _7313_/B sky130_fd_sc_hd__nor2_8
X_3799_ _7767_/Q vssd2 vssd2 vccd2 vccd2 _4312_/A sky130_fd_sc_hd__inv_2
X_5607_ _5607_/A _5607_/B vssd2 vssd2 vccd2 vccd2 _6016_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_103_137 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5538_ _5539_/A _5539_/B _5539_/C vssd2 vssd2 vccd2 vccd2 _5558_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_260 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_111_181 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7208_ _7209_/A _7209_/B vssd2 vssd2 vccd2 vccd2 _7210_/A sky130_fd_sc_hd__nand2_1
X_5469_ _5469_/A _5469_/B vssd2 vssd2 vccd2 vccd2 _5470_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__4865__B1 _5222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7139_ _7139_/A _7139_/B vssd2 vssd2 vccd2 vccd2 _7141_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_433 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1323 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1356 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_360 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_37_500 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1389 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_190 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_37_566 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xinput18 input18/A vssd2 vssd2 vccd2 vccd2 input18/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_599 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_107_487 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_91_193 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4599__A _5042_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_52_569 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xinput29 input29/A vssd2 vssd2 vccd2 vccd2 input29/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5207__B _5550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_32_293 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_671 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4320__A2 _4782_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_411 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_99_293 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_90_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_59_124 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_87_488 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_75_617 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4840_ _4841_/A _4841_/B vssd2 vssd2 vccd2 vccd2 _4842_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_511 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4771_ _4772_/A _4772_/B _4770_/Y vssd2 vssd2 vccd2 vccd2 _4920_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__5893__A _6402_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_330 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6989__A _6989_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_7_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_7_438 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_7_416 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6510_ _6510_/A _6510_/B vssd2 vssd2 vccd2 vccd2 _6510_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_55_385 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7490_ _7524_/A vssd2 vssd2 vccd2 vccd2 _7490_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_99_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6441_ _6441_/A _6441_/B vssd2 vssd2 vccd2 vccd2 _6442_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_70_355 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_43_558 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6372_ _6372_/A _6372_/B vssd2 vssd2 vccd2 vccd2 _6373_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_388 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_30_208 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_101_608 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5323_ _5324_/A _5324_/B vssd2 vssd2 vccd2 vccd2 _5388_/A sky130_fd_sc_hd__or2_1
XFILLER_0_23_293 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__7613__A _7613_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5254_ _5254_/A _5254_/B vssd2 vssd2 vccd2 vccd2 _5257_/A sky130_fd_sc_hd__xnor2_4
X_5185_ _5186_/A _5186_/B vssd2 vssd2 vccd2 vccd2 _5185_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_48_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4205_ _7765_/Q _4656_/C _4328_/B _7767_/Q _4204_/X vssd2 vssd2 vccd2 vccd2 _4206_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5133__A _5133_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4136_ _4136_/A _4136_/B vssd2 vssd2 vccd2 vccd2 _4189_/C sky130_fd_sc_hd__xor2_2
X_4067_ _4022_/B _4893_/A _4252_/C vssd2 vssd2 vccd2 vccd2 _4067_/X sky130_fd_sc_hd__and3b_1
X_7826_ _7826_/CLK _7826_/D _7585_/Y vssd2 vssd2 vccd2 vccd2 _7826_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_93_436 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_65_138 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4969_ _4969_/A _4969_/B vssd2 vssd2 vccd2 vccd2 _4970_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__5575__A1 _4893_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7757_ _7758_/CLK _7757_/D _7516_/Y vssd2 vssd2 vccd2 vccd2 _7757_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_544 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_108 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6708_ _6708_/A _6708_/B vssd2 vssd2 vccd2 vccd2 _6719_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_300 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_46_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7688_ _7800_/CLK _7688_/D vssd2 vssd2 vccd2 vccd2 _7688_/Q sky130_fd_sc_hd__dfxtp_1
X_6639_ _6039_/X _6040_/X _7143_/A _5992_/B vssd2 vssd2 vccd2 vccd2 _6641_/B sky130_fd_sc_hd__o211a_1
XANTENNA__5773__A_N _6152_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5327__A1 _4965_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_14_271 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4866__B _5210_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7523__A _7557_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout173 _4736_/A vssd2 vssd2 vccd2 vccd2 _4863_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__7252__A1 _7253_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout195 _5207_/A vssd2 vssd2 vccd2 vccd2 _5099_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__5978__A _6282_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4882__A _4882_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7252__B2 _7253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5263__B1 _4814_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_433 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1131 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_447 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XTAP_1164 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_499 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1197 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4369__A2 _4711_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_37_374 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_4_408 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_107_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4122__A _4454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_52_399 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_85_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_926 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_79_208 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6990_ _6991_/A _6991_/B vssd2 vssd2 vccd2 vccd2 _7070_/B sky130_fd_sc_hd__nand2_1
X_5941_ _7846_/Q _6357_/B _5938_/X _5939_/X _5940_/X vssd2 vssd2 vccd2 vccd2 _5947_/B
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__6215__C _6215_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_75_414 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5872_ _6071_/B _5872_/B vssd2 vssd2 vccd2 vccd2 _5883_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_0_wb_clk_i clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7795_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7611_ _7613_/A vssd2 vssd2 vccd2 vccd2 _7611_/Y sky130_fd_sc_hd__inv_2
X_4823_ _4749_/A _4749_/B _4738_/Y vssd2 vssd2 vccd2 vccd2 _4825_/B sky130_fd_sc_hd__a21bo_2
XFILLER_0_28_330 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4754_ _4673_/A _4673_/B _4671_/Y vssd2 vssd2 vccd2 vccd2 _4756_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__7608__A _7613_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_43_300 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_7_246 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7542_ _7561_/A vssd2 vssd2 vccd2 vccd2 _7542_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5309__A1 _5257_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7473_ _7713_/Q _7483_/A2 _7483_/B1 hold331/X vssd2 vssd2 vccd2 vccd2 _7473_/X sky130_fd_sc_hd__a22o_1
X_4685_ _4685_/A _4685_/B vssd2 vssd2 vccd2 vccd2 _4686_/B sky130_fd_sc_hd__or2_1
XFILLER_0_50_95 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_43_377 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6424_ _6424_/A _6424_/B _7197_/A vssd2 vssd2 vccd2 vccd2 _6426_/B sky130_fd_sc_hd__and3_1
XANTENNA__4032__A _7763_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6355_ _6668_/A _7197_/A vssd2 vssd2 vccd2 vccd2 _6365_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4389__D _5042_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5306_ _5447_/B vssd2 vssd2 vccd2 vccd2 _5308_/A sky130_fd_sc_hd__inv_2
X_6286_ _6281_/X _6284_/X _5937_/B vssd2 vssd2 vccd2 vccd2 _7237_/A sky130_fd_sc_hd__o21ai_4
X_5237_ _5183_/A _5183_/B _5181_/X vssd2 vssd2 vccd2 vccd2 _5239_/B sky130_fd_sc_hd__o21a_2
XANTENNA__5493__B1 _5550_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5168_ _5168_/A _5528_/B _5169_/B vssd2 vssd2 vccd2 vccd2 _5227_/A sky130_fd_sc_hd__or3_1
XFILLER_0_98_517 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5099_ _5099_/A _5374_/B _5100_/A vssd2 vssd2 vccd2 vccd2 _5099_/X sky130_fd_sc_hd__or3_1
X_4119_ _4882_/A _4863_/A vssd2 vssd2 vccd2 vccd2 _4132_/A sky130_fd_sc_hd__or2_1
XANTENNA__6993__B1 _6281_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_39_617 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XPHY_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_109_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XPHY_214 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_203 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_78_296 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_78_285 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_66_425 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7809_ _7814_/CLK _7809_/D _7568_/Y vssd2 vssd2 vccd2 vccd2 _7809_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_341 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7237__B _7291_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_34_322 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_104_221 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_22_528 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_104_265 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7253__A _7253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_30_572 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_55_18 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold7 hold7/A vssd2 vssd2 vccd2 vccd2 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4039__A1 _7765_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5787__A1 _5778_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_263 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5220__B _5468_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_594 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_57_425 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6035__C _6158_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_57_469 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6736__B1 _6664_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3956__A _5030_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7428__A _7436_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4211__B2 _7766_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4211__A1 _7765_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_20_43 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4470_ _4470_/A _4470_/B vssd2 vssd2 vccd2 vccd2 _4471_/B sky130_fd_sc_hd__xnor2_4
Xhold418 input29/X vssd2 vssd2 vccd2 vccd2 hold4/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6986__B _7253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold407 _7774_/Q vssd2 vssd2 vccd2 vccd2 hold407/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_54 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold429 hold5/X vssd2 vssd2 vccd2 vccd2 input2/A sky130_fd_sc_hd__dlygate4sd3_1
X_6140_ _6140_/A _6140_/B vssd2 vssd2 vccd2 vccd2 _6142_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_21_572 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_701 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_52 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_723 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _6670_/A _6071_/B vssd2 vssd2 vccd2 vccd2 _6071_/X sky130_fd_sc_hd__and2_2
XANTENNA__4278__A1 _4882_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_745 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5022_/A _5022_/B vssd2 vssd2 vccd2 vccd2 _5024_/C sky130_fd_sc_hd__xnor2_1
XTAP_789 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__6226__B _7197_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6973_ _6973_/A _6973_/B _7253_/C _7253_/D vssd2 vssd2 vccd2 vccd2 _7040_/A sky130_fd_sc_hd__or4_1
X_5924_ _6397_/A _5977_/B vssd2 vssd2 vccd2 vccd2 _5924_/X sky130_fd_sc_hd__and2_1
XFILLER_0_75_244 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6727__B1 _6430_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5855_ _5944_/C _5944_/D _5855_/C vssd2 vssd2 vccd2 vccd2 _5857_/C sky130_fd_sc_hd__and3_1
XFILLER_0_75_277 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4806_ _5164_/A _5222_/A vssd2 vssd2 vccd2 vccd2 _4808_/A sky130_fd_sc_hd__or2_2
XFILLER_0_61_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_8_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA_fanout230_A hold104/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_16_300 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__3866__A _7762_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_106_519 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_56_491 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5786_ _7846_/Q _5785_/X _5784_/X _5745_/X vssd2 vssd2 vccd2 vccd2 _5786_/Y sky130_fd_sc_hd__a211oi_4
X_4737_ _4737_/A _4737_/B vssd2 vssd2 vccd2 vccd2 _4739_/B sky130_fd_sc_hd__xnor2_1
X_7525_ _7557_/A vssd2 vssd2 vccd2 vccd2 _7525_/Y sky130_fd_sc_hd__inv_2
X_4668_ _4668_/A _4668_/B vssd2 vssd2 vccd2 vccd2 _4669_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_84 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7456_ _7696_/Q _7454_/C _7485_/B1 hold251/X vssd2 vssd2 vccd2 vccd2 _7456_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3961__B1 _4050_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6407_ _6332_/A _6329_/X _6331_/B vssd2 vssd2 vccd2 vccd2 _6409_/B sky130_fd_sc_hd__a21o_1
X_4599_ _5042_/A _5220_/A vssd2 vssd2 vccd2 vccd2 _4601_/B sky130_fd_sc_hd__nor2_1
X_7387_ _7387_/A _7420_/B _7454_/B vssd2 vssd2 vccd2 vccd2 _7387_/X sky130_fd_sc_hd__or3_1
XFILLER_0_101_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6338_ _6634_/B _6571_/B _6267_/B _6269_/A _6269_/B vssd2 vssd2 vccd2 vccd2 _6348_/A
+ sky130_fd_sc_hd__a32o_1
X_6269_ _6269_/A _6269_/B vssd2 vssd2 vccd2 vccd2 _6271_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__4269__A1 _4809_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6136__B _7037_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_79_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5040__B _5222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_109_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_81_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_62_450 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5941__A1 _7846_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_105_596 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_50_645 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4400__A _4882_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5457__B1 _4814_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6327__A _6707_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_82_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5209__B1 _5498_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_77_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4432__A1 _5042_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3970_ _4814_/B _4063_/B vssd2 vssd2 vccd2 vccd2 _3971_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_85_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4432__B2 _4863_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6709__B1 _7143_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5640_ _7858_/Q _5640_/B vssd2 vssd2 vccd2 vccd2 _6424_/A sky130_fd_sc_hd__xor2_4
XANTENNA__5932__B2 _6550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5571_ _5549_/A _5548_/B _5566_/A _5548_/A vssd2 vssd2 vccd2 vccd2 _5572_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_25_141 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_31_64 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7310_ _7310_/A _7310_/B _7310_/C vssd2 vssd2 vccd2 vccd2 _7335_/A sky130_fd_sc_hd__or3_2
XFILLER_0_25_174 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4522_ _7772_/Q _4656_/B _4522_/C vssd2 vssd2 vccd2 vccd2 _4522_/X sky130_fd_sc_hd__and3_1
X_7241_ _7242_/A _7242_/B vssd2 vssd2 vccd2 vccd2 _7275_/A sky130_fd_sc_hd__and2b_1
X_4453_ _4898_/A _5220_/A vssd2 vssd2 vccd2 vccd2 _4467_/A sky130_fd_sc_hd__or2_1
Xhold204 hold379/X vssd2 vssd2 vccd2 vccd2 _7761_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 _7427_/X vssd2 vssd2 vccd2 vccd2 _7428_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 _7449_/X vssd2 vssd2 vccd2 vccd2 _7450_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 hold612/X vssd2 vssd2 vccd2 vccd2 hold613/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 _7730_/Q vssd2 vssd2 vccd2 vccd2 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 _7457_/X vssd2 vssd2 vccd2 vccd2 _7697_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5406__A _5406_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7172_ _7211_/C _7130_/B _7126_/A vssd2 vssd2 vccd2 vccd2 _7173_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__4310__A _4898_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_21_391 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_40_188 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4384_ _4328_/A _4745_/A _4383_/X vssd2 vssd2 vccd2 vccd2 _4384_/Y sky130_fd_sc_hd__a21oi_1
X_6123_ _6184_/B _6123_/B vssd2 vssd2 vccd2 vccd2 _6311_/B sky130_fd_sc_hd__xnor2_1
XTAP_520 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6051_/X _6052_/Y _6003_/B _6003_/Y vssd2 vssd2 vccd2 vccd2 _6055_/C sky130_fd_sc_hd__o211ai_1
XANTENNA__7621__A _7627_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_553 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5005_/A _5005_/B vssd2 vssd2 vccd2 vccd2 _5005_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_56_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_586 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA_fanout278_A _7440_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5498__D _5498_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_95_317 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6956_ _6956_/A _6956_/B vssd2 vssd2 vccd2 vccd2 _6959_/A sky130_fd_sc_hd__xnor2_1
X_5907_ _6138_/A _6634_/B _6436_/A _5907_/D vssd2 vssd2 vccd2 vccd2 _5908_/A sky130_fd_sc_hd__and4b_1
XFILLER_0_91_512 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6887_ _6887_/A _6887_/B _6875_/X vssd2 vssd2 vccd2 vccd2 _6932_/A sky130_fd_sc_hd__nor3b_2
XFILLER_0_76_597 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5838_ _6283_/A _5662_/C _5920_/D _5834_/X _5837_/X vssd2 vssd2 vccd2 vccd2 _5838_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_36_439 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5769_ _6102_/B _5769_/B _6102_/C vssd2 vssd2 vccd2 vccd2 _5769_/X sky130_fd_sc_hd__and3_4
XFILLER_0_44_472 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__3934__B1 _4050_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7508_ _7565_/A vssd2 vssd2 vccd2 vccd2 _7508_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_114_393 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7439_ hold221/X _7688_/Q _7451_/S vssd2 vssd2 vccd2 vccd2 _7439_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5151__A2 _5315_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7531__A _7564_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_99_601 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6147__A _6812_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_98_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_59_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_98_177 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6403__A2 _6479_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_328 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5986__A _6092_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_67_553 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_417 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_39_277 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_82_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_82_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_22_122 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_494 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_105_393 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4130__A _4598_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_93_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4784__B _5276_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_89_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6810_ _6424_/A _6424_/B _7313_/B _7294_/C _6664_/A vssd2 vssd2 vccd2 vccd2 _6815_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_58_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4008__C _4267_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7790_ _7806_/CLK _7790_/D _7549_/Y vssd2 vssd2 vccd2 vccd2 _7790_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_309 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_85_350 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6504__B _6812_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6741_ _6741_/A _6741_/B vssd2 vssd2 vccd2 vccd2 _6742_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_586 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_45_203 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_3953_ _4050_/B _3954_/C _7779_/Q vssd2 vssd2 vccd2 vccd2 _3955_/A sky130_fd_sc_hd__a21oi_1
X_6672_ _6673_/A _6673_/B vssd2 vssd2 vccd2 vccd2 _6741_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_45_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3884_ _3864_/X _3867_/Y _3869_/X _3883_/X _7791_/Q vssd2 vssd2 vccd2 vccd2 _3904_/A
+ sky130_fd_sc_hd__o41ai_4
XFILLER_0_42_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5623_ _5618_/X _5620_/X _6071_/B _5608_/Y vssd2 vssd2 vccd2 vccd2 _5623_/X sky130_fd_sc_hd__o211a_1
XANTENNA__7616__A _7641_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_26_472 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5554_ _5528_/A _5431_/B _5553_/X vssd2 vssd2 vccd2 vccd2 _5556_/A sky130_fd_sc_hd__o21ba_1
X_4505_ _4506_/A _4506_/B vssd2 vssd2 vccd2 vccd2 _4558_/B sky130_fd_sc_hd__nand2b_1
X_5485_ _5487_/A _5487_/B vssd2 vssd2 vccd2 vccd2 _5485_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_41_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4436_ _4436_/A _4436_/B vssd2 vssd2 vccd2 vccd2 _4438_/B sky130_fd_sc_hd__xor2_4
X_7224_ _7224_/A _7255_/B vssd2 vssd2 vccd2 vccd2 _7225_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_1_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_13_188 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_111_385 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7155_ _7155_/A _7155_/B vssd2 vssd2 vccd2 vccd2 _7155_/X sky130_fd_sc_hd__or2_1
X_4367_ _4438_/A _4367_/B vssd2 vssd2 vccd2 vccd2 _4370_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_1_572 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6106_ _6106_/A _6106_/B _6106_/C vssd2 vssd2 vccd2 vccd2 _6109_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_67_71 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_350 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7086_ _7131_/A _7326_/A _7034_/A vssd2 vssd2 vccd2 vccd2 _7087_/B sky130_fd_sc_hd__a21oi_1
XTAP_394 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _4299_/A _4299_/B vssd2 vssd2 vccd2 vccd2 _4418_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6633__A2 _7253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6037_ _6100_/D _6034_/X _6035_/X _6036_/X vssd2 vssd2 vccd2 vccd2 _6037_/X sky130_fd_sc_hd__a211o_1
XTAP_1505 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_648 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_96_637 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_83_81 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_68_317 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_12 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_23 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_34 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_45 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_56 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_169 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6939_ _6939_/A _7255_/B vssd2 vssd2 vccd2 vccd2 _6940_/B sky130_fd_sc_hd__nor2_1
XPHY_89 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_67 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_78 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_76_394 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_24_409 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_17_461 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_17_472 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6430__A _6668_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6787__D _7143_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_102_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4332__B1 _4267_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold590 input44/X vssd2 vssd2 vccd2 vccd2 hold88/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_74_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4399__B1 _5099_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7337__B1 _7336_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_27_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4125__A _7767_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_103_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_82_331 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_70_504 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7436__A _7436_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6340__A _6783_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_88_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4779__B _5550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_70_548 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xoutput106 hold651/X vssd2 vssd2 vccd2 vccd2 hold292/A sky130_fd_sc_hd__buf_6
XFILLER_0_23_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xoutput117 hold663/X vssd2 vssd2 vccd2 vccd2 hold310/A sky130_fd_sc_hd__buf_6
Xoutput128 hold619/X vssd2 vssd2 vccd2 vccd2 hold266/A sky130_fd_sc_hd__buf_6
X_5270_ _5270_/A _5270_/B vssd2 vssd2 vccd2 vccd2 _5272_/B sky130_fd_sc_hd__xor2_1
Xoutput139 _7709_/Q vssd2 vssd2 vccd2 vccd2 wbs_dat_o[14] sky130_fd_sc_hd__buf_12
XANTENNA__6863__A2 _7145_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4221_ _4221_/A _4221_/B vssd2 vssd2 vccd2 vccd2 _4234_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_41 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4152_ _7766_/Q _4454_/B vssd2 vssd2 vccd2 vccd2 _4152_/X sky130_fd_sc_hd__and2_1
XFILLER_0_37_63 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4083_ _7763_/Q _4083_/B _4146_/B vssd2 vssd2 vccd2 vccd2 _4083_/X sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_96 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7842_ _7854_/CLK _7842_/D _7601_/Y vssd2 vssd2 vccd2 vccd2 _7842_/Q sky130_fd_sc_hd__dfrtp_4
X_4985_ _4985_/A _4985_/B vssd2 vssd2 vccd2 vccd2 _4986_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_77_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7773_ _7804_/CLK _7773_/D _7532_/Y vssd2 vssd2 vccd2 vccd2 _7773_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6724_ _6724_/A _6724_/B vssd2 vssd2 vccd2 vccd2 _6750_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_512 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3936_ _7783_/Q _3936_/B vssd2 vssd2 vccd2 vccd2 _4162_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_73_353 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_73_397 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6655_ _6973_/A _6973_/B _7045_/A _7140_/A vssd2 vssd2 vccd2 vccd2 _6656_/B sky130_fd_sc_hd__or4_1
XFILLER_0_46_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3867_ _3865_/Y _3866_/Y _4656_/C vssd2 vssd2 vccd2 vccd2 _3867_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6586_ _5816_/A _5816_/B _7253_/C vssd2 vssd2 vccd2 vccd2 _6591_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_33_239 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_3798_ _7768_/Q vssd2 vssd2 vccd2 vccd2 _4374_/A sky130_fd_sc_hd__inv_2
X_5606_ _7866_/Q _5612_/B _5606_/C vssd2 vssd2 vccd2 vccd2 _5828_/C sky130_fd_sc_hd__or3_4
XFILLER_0_14_464 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5537_ _5537_/A _5537_/B vssd2 vssd2 vccd2 vccd2 _5539_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_103_149 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_41_272 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7207_ _7168_/A _7168_/B _7167_/A vssd2 vssd2 vccd2 vccd2 _7209_/B sky130_fd_sc_hd__a21o_1
X_5468_ _5468_/A _5550_/A vssd2 vssd2 vccd2 vccd2 _5469_/B sky130_fd_sc_hd__or2_1
XFILLER_0_111_193 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4865__A1 _5210_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4865__B2 _5210_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5399_ _5401_/A vssd2 vssd2 vccd2 vccd2 _5445_/B sky130_fd_sc_hd__inv_2
X_4419_ _4419_/A vssd2 vssd2 vccd2 vccd2 _4420_/B sky130_fd_sc_hd__inv_2
X_7138_ _7237_/A _7224_/A _7138_/C _7253_/B vssd2 vssd2 vccd2 vccd2 _7139_/B sky130_fd_sc_hd__or4_1
X_7069_ _7070_/A _7070_/B _7070_/C vssd2 vssd2 vccd2 vccd2 _7123_/A sky130_fd_sc_hd__a21oi_2
XTAP_1313 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6425__A _6425_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_68_136 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_96_489 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_96_467 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1357 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1379 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_353 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_107_455 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_107_444 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_91_161 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
Xinput19 input19/A vssd2 vssd2 vccd2 vccd2 input19/X sky130_fd_sc_hd__buf_1
XANTENNA__4599__B _5220_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_52_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_32_283 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_99_261 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_90_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_59_136 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_59_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_23_10 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_23_21 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_74_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_23_43 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_28_523 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4770_ _4709_/A _4709_/B _4705_/B vssd2 vssd2 vccd2 vccd2 _4770_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__5893__B _6150_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_342 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__6989__B _7255_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_70_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_99_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6440_ _6441_/A _6441_/B vssd2 vssd2 vccd2 vccd2 _6440_/X sky130_fd_sc_hd__and2_1
XFILLER_0_82_194 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_55_397 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_43_548 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_113_447 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6371_ _6372_/A _6372_/B vssd2 vssd2 vccd2 vccd2 _6371_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_51_570 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5322_ _5281_/A _5281_/B _5288_/Y vssd2 vssd2 vccd2 vccd2 _5324_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_11_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5253_ _4996_/B _5249_/X _5252_/Y vssd2 vssd2 vccd2 vccd2 _5254_/B sky130_fd_sc_hd__a21o_2
X_5184_ _5115_/A _5115_/B _5113_/X vssd2 vssd2 vccd2 vccd2 _5186_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_48_62 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__5414__A _5414_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4204_ _7766_/Q _4745_/A _5458_/A vssd2 vssd2 vccd2 vccd2 _4204_/X sky130_fd_sc_hd__and3_1
X_4135_ _4135_/A _4135_/B vssd2 vssd2 vccd2 vccd2 _4136_/B sky130_fd_sc_hd__nand2_1
X_4066_ _4268_/A _4122_/D _4066_/C _4066_/D vssd2 vssd2 vccd2 vccd2 _4066_/X sky130_fd_sc_hd__and4_1
X_7825_ _7826_/CLK _7825_/D _7584_/Y vssd2 vssd2 vccd2 vccd2 _7825_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4061__D_N _7766_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_38_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_93_426 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_59_670 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_19_512 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_19_523 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4968_ _4969_/A _4969_/B vssd2 vssd2 vccd2 vccd2 _4968_/Y sky130_fd_sc_hd__nand2_1
X_7756_ _7758_/CLK _7756_/D _7515_/Y vssd2 vssd2 vccd2 vccd2 _7756_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5575__A2 _4006_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6707_ _6707_/A _7255_/B vssd2 vssd2 vccd2 vccd2 _6708_/B sky130_fd_sc_hd__nor2_1
X_4899_ _4899_/A _4899_/B vssd2 vssd2 vccd2 vccd2 _4900_/B sky130_fd_sc_hd__xnor2_4
X_7687_ _7782_/CLK _7687_/D vssd2 vssd2 vccd2 vccd2 _7687_/Q sky130_fd_sc_hd__dfxtp_1
X_3919_ _4252_/B _4252_/C _7764_/Q vssd2 vssd2 vccd2 vccd2 _3919_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_61_345 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6638_ _5991_/X _5993_/X _7143_/B _5781_/B vssd2 vssd2 vccd2 vccd2 _6641_/A sky130_fd_sc_hd__o211a_1
XFILLER_0_34_537 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5327__A2 _5528_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6569_ _6505_/A _6507_/B _6505_/B vssd2 vssd2 vccd2 vccd2 _6574_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__4866__C _4965_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout174 _4779_/A vssd2 vssd2 vccd2 vccd2 _4898_/A sky130_fd_sc_hd__buf_4
Xfanout196 _4318_/Y vssd2 vssd2 vccd2 vccd2 _4782_/B sky130_fd_sc_hd__buf_4
XFILLER_0_88_209 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7252__A2 _7253_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_96_253 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1132 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_489 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1198 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_673 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_37_353 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_654 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_52_334 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_37_386 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_69_28 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_40_507 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_20_220 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_916 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_264 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_85_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_949 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_9 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5940_ _7845_/Q _6283_/B _6587_/B vssd2 vssd2 vccd2 vccd2 _5940_/X sky130_fd_sc_hd__and3_1
XANTENNA__6215__D _6989_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7610_ _7613_/A vssd2 vssd2 vccd2 vccd2 _7610_/Y sky130_fd_sc_hd__inv_2
X_5871_ _6670_/A _6019_/D _5834_/B _7846_/Q _6016_/B vssd2 vssd2 vccd2 vccd2 _5872_/B
+ sky130_fd_sc_hd__a32o_1
X_4822_ _4822_/A _4822_/B vssd2 vssd2 vccd2 vccd2 _4825_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_90_429 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4753_ _4753_/A _4753_/B vssd2 vssd2 vccd2 vccd2 _4756_/A sky130_fd_sc_hd__xnor2_1
X_7541_ _7561_/A vssd2 vssd2 vccd2 vccd2 _7541_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_504 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_16_515 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7472_ _7712_/Q _7483_/A2 _7483_/B1 hold335/X vssd2 vssd2 vccd2 vccd2 _7472_/X sky130_fd_sc_hd__a22o_1
X_6423_ _6425_/A _7094_/A vssd2 vssd2 vccd2 vccd2 _6426_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_665 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4684_ _4685_/A _4685_/B vssd2 vssd2 vccd2 vccd2 _4686_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__7624__A _7627_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6354_ _6354_/A _6354_/B vssd2 vssd2 vccd2 vccd2 _6369_/A sky130_fd_sc_hd__xor2_2
X_5305_ _5305_/A _5305_/B vssd2 vssd2 vccd2 vccd2 _5447_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__3871__B _5458_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6285_ _6281_/X _6284_/X _5937_/B vssd2 vssd2 vccd2 vccd2 _6430_/B sky130_fd_sc_hd__o21a_4
XANTENNA__5144__A _5145_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5236_ _5295_/B _5236_/B vssd2 vssd2 vccd2 vccd2 _5239_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_52_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7482__A2 _7483_/A2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5493__A1 _5468_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5167_ _4380_/Y _4382_/X _4385_/X _5374_/B _4144_/D vssd2 vssd2 vccd2 vccd2 _5169_/B
+ sky130_fd_sc_hd__a311o_1
X_5098_ _4327_/X _4331_/X _5326_/B _4267_/D vssd2 vssd2 vccd2 vccd2 _5100_/B sky130_fd_sc_hd__o211a_1
X_4118_ _4118_/A _4118_/B vssd2 vssd2 vccd2 vccd2 _4136_/A sky130_fd_sc_hd__xnor2_2
X_4049_ _7806_/Q _4049_/B vssd2 vssd2 vccd2 vccd2 _4049_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_66_404 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_215 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_204 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_93_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_91_81 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_226 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7808_ _7814_/CLK _7808_/D _7567_/Y vssd2 vssd2 vccd2 vccd2 _7808_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_109 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7739_ _7739_/CLK _7739_/D _7498_/Y vssd2 vssd2 vccd2 vccd2 _7739_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_194 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_34_334 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_62_665 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_104_233 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_61_186 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__7534__A _7557_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_15_570 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_34_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_104_277 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7253__B _7253_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7473__A2 _7483_/A2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4893__A _4893_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold8 hold8/A vssd2 vssd2 vccd2 vccd2 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_518 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_69_220 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_97_540 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5787__A2 _5786_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_29_117 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_84_256 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_44_109 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_65_492 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_80_451 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_53_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_53_665 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_20_11 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_20_33 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_111_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_80_473 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xhold408 wbs_dat_i[9] vssd2 vssd2 vccd2 vccd2 hold408/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold419 hold4/X vssd2 vssd2 vccd2 vccd2 _7842_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7444__A _7452_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_21_551 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_702 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6029_/A _6029_/B _6031_/X vssd2 vssd2 vccd2 vccd2 _6086_/A sky130_fd_sc_hd__a21bo_1
XTAP_768 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7464__A2 _7454_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_29_75 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4278__A2 _4896_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_735 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5021_/A _5021_/B vssd2 vssd2 vccd2 vccd2 _5022_/B sky130_fd_sc_hd__xor2_1
XTAP_779 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6972_ _6571_/B _7294_/C _7313_/B _6571_/A vssd2 vssd2 vccd2 vccd2 _6974_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_88_573 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_48_426 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5923_ _5923_/A _5923_/B _5923_/C _5923_/D vssd2 vssd2 vccd2 vccd2 _5923_/X sky130_fd_sc_hd__or4_1
XFILLER_0_61_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6727__A1 _6571_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6727__B2 _6571_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_48_448 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5854_ _5845_/X _5846_/Y _5944_/C vssd2 vssd2 vccd2 vccd2 _5857_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_75_267 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4805_ _4805_/A _4805_/B vssd2 vssd2 vccd2 vccd2 _4826_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_61_62 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7524_ _7524_/A vssd2 vssd2 vccd2 vccd2 _7524_/Y sky130_fd_sc_hd__inv_2
X_5785_ _6152_/B _6152_/C _6281_/C vssd2 vssd2 vccd2 vccd2 _5785_/X sky130_fd_sc_hd__and3_4
XANTENNA__5950__A2 _6634_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4736_ _4736_/A _5374_/B _4737_/B vssd2 vssd2 vccd2 vccd2 _4821_/A sky130_fd_sc_hd__or3_2
XANTENNA_fanout223_A _4460_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4667_ _4896_/A _5220_/A _4668_/A vssd2 vssd2 vccd2 vccd2 _4739_/A sky130_fd_sc_hd__or3_1
XFILLER_0_43_164 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7455_ _7695_/Q _7454_/C _7485_/B1 hold249/X vssd2 vssd2 vccd2 vccd2 _7455_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3882__A _7767_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_31_326 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6406_ _6406_/A _6406_/B vssd2 vssd2 vccd2 vccd2 _6409_/A sky130_fd_sc_hd__xnor2_4
X_7386_ _7386_/A hold99/X vssd2 vssd2 vccd2 vccd2 _7386_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_540 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7354__A _7436_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6337_ _6337_/A _6337_/B vssd2 vssd2 vccd2 vccd2 _6377_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_101_225 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4598_ _4598_/A _5374_/B vssd2 vssd2 vccd2 vccd2 _4601_/A sky130_fd_sc_hd__nor2_1
X_6268_ _6707_/A _7037_/A vssd2 vssd2 vccd2 vccd2 _6269_/B sky130_fd_sc_hd__nor2_1
XANTENNA__7455__A2 _7454_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6199_ _6199_/A _6199_/B _6199_/C vssd2 vssd2 vccd2 vccd2 _6200_/B sky130_fd_sc_hd__nor3_1
X_5219_ _5219_/A _5219_/B vssd2 vssd2 vccd2 vccd2 _5235_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__5602__A _5645_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6415__B1 _6973_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_94_576 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_47_492 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6152__B _6152_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_62_484 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_34_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__3792__A _4893_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4400__B _5099_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6654__B1 _7197_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6327__B _6479_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5209__B2 _5210_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5209__A1 _5210_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_15_44 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_97_381 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__4432__A2 _4711_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6709__A1 _6039_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_15_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_85_587 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_45_407 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_110_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5932__A2 _6812_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5570_ _5570_/A _5570_/B _5570_/C vssd2 vssd2 vccd2 vccd2 _5572_/A sky130_fd_sc_hd__or3_1
XFILLER_0_31_54 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4798__A _4882_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_53_462 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_25_153 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4521_ _4521_/A _4656_/B vssd2 vssd2 vccd2 vccd2 _4521_/Y sky130_fd_sc_hd__nor2_1
X_7240_ _7270_/A _7240_/B vssd2 vssd2 vccd2 vccd2 _7242_/B sky130_fd_sc_hd__and2_1
X_4452_ _4452_/A _4452_/B vssd2 vssd2 vccd2 vccd2 _4469_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_53_495 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_13_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold216 hold401/X vssd2 vssd2 vccd2 vccd2 _7773_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 _7357_/X vssd2 vssd2 vccd2 vccd2 _7358_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_112 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold227 hold355/X vssd2 vssd2 vccd2 vccd2 _7784_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 _7458_/X vssd2 vssd2 vccd2 vccd2 _7698_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 _7727_/Q vssd2 vssd2 vccd2 vccd2 hold249/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5406__B _5550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_40_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7171_ _7214_/B _7171_/B vssd2 vssd2 vccd2 vccd2 _7211_/D sky130_fd_sc_hd__nand2_2
XANTENNA__4310__B _4711_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4383_ _7770_/Q _4656_/B _4522_/C vssd2 vssd2 vccd2 vccd2 _4383_/X sky130_fd_sc_hd__and3_1
X_6122_ _6128_/A _6122_/B vssd2 vssd2 vccd2 vccd2 _6123_/B sky130_fd_sc_hd__nor2_1
XTAP_510 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6003_/B _6003_/Y _6051_/X _6052_/Y vssd2 vssd2 vccd2 vccd2 _6055_/B sky130_fd_sc_hd__a211o_1
XTAP_554 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _5005_/A _5005_/B vssd2 vssd2 vccd2 vccd2 _5123_/A sky130_fd_sc_hd__or2_4
XTAP_587 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout173_A _4736_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_95_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6955_ _6956_/A _6956_/B vssd2 vssd2 vccd2 vccd2 _7007_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_76_543 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_76_521 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5906_ _6105_/B _6707_/A _6634_/B _6436_/A vssd2 vssd2 vccd2 vccd2 _5909_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__6253__A _6253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_76_587 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_76_565 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6886_ _6885_/B _6885_/C _6885_/A vssd2 vssd2 vccd2 vccd2 _6887_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_237 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_17_610 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_29_492 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5837_ _6253_/B _6253_/C _5827_/X _5825_/X _6157_/A vssd2 vssd2 vccd2 vccd2 _5837_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_91_557 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5768_ _6105_/A _6550_/A vssd2 vssd2 vccd2 vccd2 _7807_/D sky130_fd_sc_hd__nor2_2
XANTENNA__4204__C _5458_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4719_ _4720_/A _4720_/B vssd2 vssd2 vccd2 vccd2 _4772_/A sky130_fd_sc_hd__and2_1
X_7507_ _7565_/A vssd2 vssd2 vccd2 vccd2 _7507_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_31_101 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_114_361 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_71_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7438_ _7440_/A _7438_/B vssd2 vssd2 vccd2 vccd2 _7687_/D sky130_fd_sc_hd__and2_1
X_5699_ _7883_/Q _5699_/B vssd2 vssd2 vccd2 vccd2 _6094_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_16_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_102_523 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7369_ hold121/X _7767_/D _7383_/S vssd2 vssd2 vccd2 vccd2 _7369_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6147__B _6812_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_98_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_86_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5986__B _6783_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_79_370 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_39_234 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_109_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_54_204 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_429 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_35_440 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_35_462 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_112_309 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_105_361 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_62_292 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4130__B _5029_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_93_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_89_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6740_ _6668_/A _7313_/B _6669_/X _5907_/D vssd2 vssd2 vccd2 vccd2 _6741_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_85_362 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__6504__C _7140_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_58_554 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3952_ _7780_/Q _3952_/B vssd2 vssd2 vccd2 vccd2 _4164_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_42_42 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_73_513 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6671_ _5907_/D _7313_/B _6669_/X _6590_/A vssd2 vssd2 vccd2 vccd2 _6673_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_58_598 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3883_ _3880_/X _3881_/X _3882_/X _4326_/D vssd2 vssd2 vccd2 vccd2 _3883_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_73_579 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5622_ _5586_/B _5584_/Y _5586_/Y _5599_/B _5653_/C vssd2 vssd2 vccd2 vccd2 _6071_/B
+ sky130_fd_sc_hd__o2111a_4
XANTENNA__4169__B2 _7766_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4169__A1 _7764_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_60_218 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5553_ _5553_/A _5553_/B vssd2 vssd2 vccd2 vccd2 _5553_/X sky130_fd_sc_hd__xor2_1
X_4504_ _4504_/A _4504_/B vssd2 vssd2 vccd2 vccd2 _4506_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5484_ _5486_/A _5486_/B vssd2 vssd2 vccd2 vccd2 _5487_/B sky130_fd_sc_hd__nand2_1
X_4435_ _4435_/A _4435_/B vssd2 vssd2 vccd2 vccd2 _4436_/B sky130_fd_sc_hd__nor2_2
X_7223_ _7223_/A _7223_/B vssd2 vssd2 vccd2 vccd2 _7225_/A sky130_fd_sc_hd__nor2_1
X_7154_ _7155_/A _7155_/B vssd2 vssd2 vccd2 vccd2 _7154_/Y sky130_fd_sc_hd__nand2_1
X_4366_ _4898_/A _4863_/A _4711_/A _4782_/B vssd2 vssd2 vccd2 vccd2 _4438_/A sky130_fd_sc_hd__or4_4
XANTENNA__7632__A _7641_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6105_ _6105_/A _6105_/B _6989_/A _7047_/A vssd2 vssd2 vccd2 vccd2 _6106_/C sky130_fd_sc_hd__or4b_1
XTAP_351 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_97 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7085_ _7131_/B _7131_/C vssd2 vssd2 vccd2 vccd2 _7087_/A sky130_fd_sc_hd__and2_1
XANTENNA__5152__A _5276_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_384 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _4297_/A _4363_/A vssd2 vssd2 vccd2 vccd2 _4299_/B sky130_fd_sc_hd__xnor2_2
XTAP_395 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _7847_/Q _6283_/B vssd2 vssd2 vccd2 vccd2 _6036_/X sky130_fd_sc_hd__and2_1
XTAP_1506 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XPHY_13 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_137 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XPHY_24 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_35 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_46 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_76_362 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6938_ _6938_/A _6938_/B vssd2 vssd2 vccd2 vccd2 _6940_/A sky130_fd_sc_hd__xor2_2
XPHY_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_68 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_79 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_76_373 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_64_513 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6869_ _6916_/A _6869_/B vssd2 vssd2 vccd2 vccd2 _6871_/B sky130_fd_sc_hd__or2_1
XANTENNA__6711__A _6989_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_36_237 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_91_376 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_51_229 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6430__B _6430_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_44_292 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_32_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6857__B1 _7143_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold580 la_data_in[33] vssd2 vssd2 vccd2 vccd2 hold77/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6872__A3 _6669_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold591 hold88/X vssd2 vssd2 vccd2 vccd2 _7876_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6158__A _6158_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5832__B2 _7844_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5832__A1 _7842_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_649 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_86_126 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_95_671 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_67_373 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__7337__B2 _7336_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_568 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_12_23 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_237 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_103_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_70_516 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_12_67 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5899__B2 _6158_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5899__A1 _7847_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6340__B _7037_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_88_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_42_229 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_112_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xoutput107 hold647/X vssd2 vssd2 vccd2 vccd2 hold298/A sky130_fd_sc_hd__buf_6
Xoutput118 hold665/X vssd2 vssd2 vccd2 vccd2 hold312/A sky130_fd_sc_hd__buf_6
Xoutput129 hold613/X vssd2 vssd2 vccd2 vccd2 hold260/A sky130_fd_sc_hd__buf_6
XFILLER_0_11_627 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7452__A _7452_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4220_ _4220_/A _4220_/B vssd2 vssd2 vccd2 vccd2 _4221_/B sky130_fd_sc_hd__and2_1
X_4151_ _4142_/X _4145_/X _4149_/X _3880_/A vssd2 vssd2 vccd2 vccd2 _4155_/B sky130_fd_sc_hd__a31o_1
X_4082_ _4656_/A _4082_/B _4083_/B _4082_/D vssd2 vssd2 vccd2 vccd2 _4082_/X sky130_fd_sc_hd__and4_1
XFILLER_0_37_53 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_37_75 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7841_ _7854_/CLK _7841_/D _7600_/Y vssd2 vssd2 vccd2 vccd2 _7841_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_53_52 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4984_ _4985_/A _4985_/B vssd2 vssd2 vccd2 vccd2 _4984_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_77_159 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7772_ _7806_/CLK _7772_/D _7531_/Y vssd2 vssd2 vccd2 vccd2 _7772_/Q sky130_fd_sc_hd__dfrtp_4
X_6723_ _6724_/A _6724_/B vssd2 vssd2 vccd2 vccd2 _6776_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_73_310 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_58_373 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_46_524 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3935_ _7784_/Q _3935_/B vssd2 vssd2 vccd2 vccd2 _4022_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_85_181 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6654_ _6571_/B _7094_/A _7197_/A _6571_/A vssd2 vssd2 vccd2 vccd2 _6656_/A sky130_fd_sc_hd__a22o_1
XANTENNA__7627__A _7627_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_61_505 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_3866_ _7762_/Q _4656_/B _4454_/B vssd2 vssd2 vccd2 vccd2 _3866_/Y sky130_fd_sc_hd__nand3_1
X_5605_ _7866_/Q _5612_/B _5606_/C vssd2 vssd2 vccd2 vccd2 _5607_/B sky130_fd_sc_hd__nor3_2
XFILLER_0_82_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6585_ _6668_/A _7222_/B vssd2 vssd2 vccd2 vccd2 _6592_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_549 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_538 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3797_ _4328_/A vssd2 vssd2 vccd2 vccd2 _4149_/A sky130_fd_sc_hd__inv_2
XFILLER_0_14_454 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5536_ _5468_/A _5431_/B _5499_/B vssd2 vssd2 vccd2 vccd2 _5537_/B sky130_fd_sc_hd__o21ai_1
X_5467_ _5498_/A _5528_/A _5550_/B _5404_/A vssd2 vssd2 vccd2 vccd2 _5469_/A sky130_fd_sc_hd__o22a_1
XFILLER_0_111_161 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7206_ _7246_/B _7206_/B vssd2 vssd2 vccd2 vccd2 _7209_/A sky130_fd_sc_hd__nor2_1
XANTENNA__7362__A _7440_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4418_ _4418_/A _4418_/B vssd2 vssd2 vccd2 vccd2 _4419_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_41_295 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4865__A2 _4965_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5398_ _5398_/A _5398_/B vssd2 vssd2 vccd2 vccd2 _5401_/A sky130_fd_sc_hd__xor2_4
X_7137_ _7099_/B _7222_/A _7222_/C _6430_/B vssd2 vssd2 vccd2 vccd2 _7139_/A sky130_fd_sc_hd__a22o_1
X_4349_ _4350_/A _4350_/B vssd2 vssd2 vccd2 vccd2 _4408_/A sky130_fd_sc_hd__nand2_1
X_7068_ _7004_/A _7004_/B _7002_/X vssd2 vssd2 vccd2 vccd2 _7070_/C sky130_fd_sc_hd__a21oi_2
X_6019_ _6398_/A _6071_/B _6019_/C _6019_/D vssd2 vssd2 vccd2 vccd2 _6019_/X sky130_fd_sc_hd__and4_1
XTAP_1314 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6425__B _7094_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1347 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_470 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_37_557 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_64_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_52_549 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_17_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_60_593 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_58_19 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4896__A _4896_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_20_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_74_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_99_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_87_457 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_59_148 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_114_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6230__A1 _6668_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_28_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_99_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6351__A _6812_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_43_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_70_324 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6370_ _6295_/A _6293_/Y _6292_/Y vssd2 vssd2 vccd2 vccd2 _6372_/B sky130_fd_sc_hd__o21ai_2
X_5321_ _5370_/B _5321_/B vssd2 vssd2 vccd2 vccd2 _5324_/A sky130_fd_sc_hd__or2_1
XFILLER_0_100_109 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5252_ _5252_/A _5252_/B vssd2 vssd2 vccd2 vccd2 _5252_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_11_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5183_ _5183_/A _5183_/B vssd2 vssd2 vccd2 vccd2 _5186_/A sky130_fd_sc_hd__xnor2_2
X_4203_ _4328_/A _4458_/D _4268_/D vssd2 vssd2 vccd2 vccd2 _4206_/C sky130_fd_sc_hd__and3_1
XANTENNA__5133__C _5133_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4134_ _4134_/A _4134_/B vssd2 vssd2 vccd2 vccd2 _4135_/B sky130_fd_sc_hd__or2_1
X_4065_ _4062_/Y _4064_/X _4814_/B vssd2 vssd2 vccd2 vccd2 _4065_/X sky130_fd_sc_hd__o21a_1
X_7824_ _7826_/CLK _7824_/D _7583_/Y vssd2 vssd2 vccd2 vccd2 _7824_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_457 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_66_608 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4046__A _4598_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_fanout253_A _7886_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6221__B2 _7850_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6221__A1 _6158_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_108_209 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_93_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4967_ _4088_/A _4088_/B _5528_/B vssd2 vssd2 vccd2 vccd2 _4969_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_46_321 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7755_ _7758_/CLK _7755_/D _7514_/Y vssd2 vssd2 vccd2 vccd2 _7755_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_162 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6706_ _6704_/X _6706_/B vssd2 vssd2 vccd2 vccd2 _6708_/A sky130_fd_sc_hd__and2b_1
X_4898_ _4898_/A _5528_/B _4899_/A vssd2 vssd2 vccd2 vccd2 _4898_/X sky130_fd_sc_hd__or3_1
XFILLER_0_46_354 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7686_ _7798_/CLK _7686_/D vssd2 vssd2 vccd2 vccd2 _7686_/Q sky130_fd_sc_hd__dfxtp_1
X_3918_ _7785_/Q _3918_/B vssd2 vssd2 vccd2 vccd2 _4252_/C sky130_fd_sc_hd__xnor2_2
X_6637_ _6637_/A _6637_/B vssd2 vssd2 vccd2 vccd2 _6647_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_324 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3849_ _7792_/Q _7791_/Q _3888_/B vssd2 vssd2 vccd2 vccd2 _3851_/B sky130_fd_sc_hd__o21a_2
X_6568_ _6939_/A _6572_/B _6498_/A _6495_/X vssd2 vssd2 vccd2 vccd2 _6576_/A sky130_fd_sc_hd__o31a_1
XFILLER_0_104_448 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_89_81 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_14_262 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5519_ _5451_/A _5451_/B _5518_/Y vssd2 vssd2 vccd2 vccd2 _5561_/B sky130_fd_sc_hd__a21o_1
X_6499_ _6500_/A _6500_/B _6500_/C vssd2 vssd2 vccd2 vccd2 _6499_/X sky130_fd_sc_hd__o21a_1
XANTENNA__7092__A _7140_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_100_632 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7485__B1 _7485_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_100_654 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4866__D _5222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout175 _4747_/A vssd2 vssd2 vccd2 vccd2 _4810_/A sky130_fd_sc_hd__buf_4
Xfanout186 _6425_/A vssd2 vssd2 vccd2 vccd2 _6664_/A sky130_fd_sc_hd__clkbuf_8
Xfanout197 _4318_/Y vssd2 vssd2 vccd2 vccd2 _5210_/B sky130_fd_sc_hd__buf_4
XFILLER_0_96_221 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1111 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_479 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_96_265 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1155 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_192 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__3795__A _7771_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_37_332 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_92_460 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_25_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_37_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_92_493 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_64_184 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_52_368 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_100_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_917 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7476__B1 _7483_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_20_243 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_85_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_939 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_57 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4462__B1 _5099_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5870_ _7336_/A _5866_/Y _5867_/X _5918_/A vssd2 vssd2 vccd2 vccd2 _7809_/D sky130_fd_sc_hd__o22ai_1
XFILLER_0_75_427 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4821_ _4821_/A _4821_/B vssd2 vssd2 vccd2 vccd2 _4822_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_75_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6081__A _6550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_90_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4752_ _4752_/A _4752_/B vssd2 vssd2 vccd2 vccd2 _4753_/B sky130_fd_sc_hd__xor2_1
X_7540_ _7561_/A vssd2 vssd2 vccd2 vccd2 _7540_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_28_376 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4683_ _4683_/A _4683_/B vssd2 vssd2 vccd2 vccd2 _4685_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_173 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_43_313 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7471_ _7711_/Q _7483_/A2 _7483_/B1 hold329/X vssd2 vssd2 vccd2 vccd2 _7471_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_16_538 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6422_ _6422_/A _6422_/B vssd2 vssd2 vccd2 vccd2 _6446_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_154 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_113_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_31_519 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6353_ _6353_/A _6353_/B vssd2 vssd2 vccd2 vccd2 _6354_/B sky130_fd_sc_hd__xnor2_2
X_5304_ _5305_/A _5305_/B vssd2 vssd2 vccd2 vccd2 _5304_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_73 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7467__B1 _7485_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6284_ _6093_/A _6357_/B _5853_/C _6282_/X _6283_/X vssd2 vssd2 vccd2 vccd2 _6284_/X
+ sky130_fd_sc_hd__a2111o_2
XANTENNA__5144__B _5145_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5235_ _5235_/A _5235_/B vssd2 vssd2 vccd2 vccd2 _5236_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_45_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7640__A _7641_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5493__A2 _5528_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_75_61 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5166_ _4199_/X _4200_/X _4206_/X _4814_/Y _4080_/D vssd2 vssd2 vccd2 vccd2 _5169_/A
+ sky130_fd_sc_hd__o311a_1
XANTENNA__6256__A _7143_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4117_ _4118_/A _4118_/B vssd2 vssd2 vccd2 vccd2 _4180_/A sky130_fd_sc_hd__nand2_1
X_5097_ _4155_/A _4155_/B _4155_/C _5528_/B vssd2 vssd2 vccd2 vccd2 _5100_/A sky130_fd_sc_hd__a31o_1
X_4048_ _4053_/B _4048_/B vssd2 vssd2 vccd2 vccd2 _4052_/A sky130_fd_sc_hd__nand2_1
XPHY_216 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_205 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_91_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_78_265 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_66_416 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XPHY_227 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5999_ _5998_/B _5998_/C _5998_/A vssd2 vssd2 vccd2 vccd2 _6001_/B sky130_fd_sc_hd__a21o_1
X_7807_ _7814_/CLK _7807_/D _7566_/Y vssd2 vssd2 vccd2 vccd2 _7807_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7738_ _7739_/CLK _7738_/D _7497_/Y vssd2 vssd2 vccd2 vccd2 _7738_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4223__B _4898_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4508__A1 _4810_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_61_143 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_121 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7669_ _7782_/CLK _7669_/D vssd2 vssd2 vccd2 vccd2 _7669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_508 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_104_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_104_289 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7253__C _7253_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7458__B1 _7485_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_30_563 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7550__A _7557_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold9 hold9/A vssd2 vssd2 vccd2 vccd2 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4692__B1 _5455_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6433__A1 _6253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_276 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_57_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_37_140 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_108_540 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_13_508 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_25_357 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_111_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_80_485 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
Xhold409 _7806_/Q vssd2 vssd2 vccd2 vccd2 _4050_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_379 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_40_305 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_33_390 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_96_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_703 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5021_/A _5021_/B vssd2 vssd2 vccd2 vccd2 _5020_/Y sky130_fd_sc_hd__nor2_1
XTAP_758 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6076__A _6093_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_88_552 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_88_541 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6971_ _6571_/B _7222_/B _6922_/B _6924_/Y vssd2 vssd2 vccd2 vccd2 _6979_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_88_585 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_48_405 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__4027__C _5030_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5922_ _6282_/A _6253_/C _6075_/C _6075_/D vssd2 vssd2 vccd2 vccd2 _5923_/D sky130_fd_sc_hd__and4_1
XANTENNA__6727__A2 _7197_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5853_ _5853_/A _5853_/B _5853_/C vssd2 vssd2 vccd2 vccd2 _5853_/X sky130_fd_sc_hd__and3_1
X_4804_ _4804_/A _4804_/B vssd2 vssd2 vccd2 vccd2 _4805_/B sky130_fd_sc_hd__or2_2
X_5784_ _7844_/Q _5780_/X _5782_/X _5783_/X _5779_/X vssd2 vssd2 vccd2 vccd2 _5784_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_61_96 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4735_ _4966_/A _5220_/A vssd2 vssd2 vccd2 vccd2 _4737_/B sky130_fd_sc_hd__or2_1
X_7523_ _7557_/A vssd2 vssd2 vccd2 vccd2 _7523_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7635__A _7641_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_28_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4666_ _4896_/A _5220_/A vssd2 vssd2 vccd2 vccd2 _4668_/B sky130_fd_sc_hd__nor2_1
X_7454_ _7454_/A _7454_/B _7454_/C vssd2 vssd2 vccd2 vccd2 _7454_/Y sky130_fd_sc_hd__nor3_2
X_6405_ _6405_/A _6405_/B vssd2 vssd2 vccd2 vccd2 _6406_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_43_198 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7385_ _7349_/A _7385_/B vssd2 vssd2 vccd2 vccd2 _7385_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__6360__B1 _6281_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4597_ _4594_/X _4595_/X _4252_/B vssd2 vssd2 vccd2 vccd2 _5414_/B sky130_fd_sc_hd__o21ai_2
X_6336_ _6337_/A _6337_/B vssd2 vssd2 vccd2 vccd2 _6453_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_101_237 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6267_ _6267_/A _6267_/B vssd2 vssd2 vccd2 vccd2 _6269_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__7370__A _7452_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6198_ _6199_/A _6199_/B _6199_/C vssd2 vssd2 vccd2 vccd2 _6307_/A sky130_fd_sc_hd__o21a_1
X_5218_ _5219_/B _5219_/A vssd2 vssd2 vccd2 vccd2 _5260_/A sky130_fd_sc_hd__nand2b_1
X_5149_ _5149_/A _5149_/B vssd2 vssd2 vccd2 vccd2 _5154_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__6415__B2 _6939_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6415__A1 _6973_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_94_555 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_94_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_66_224 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_109_337 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_105_576 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_105_565 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_62_496 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_30_360 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6654__A1 _6571_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6654__B2 _6571_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4665__B1 _5374_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_89_305 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_82_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5209__A2 _5528_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6811__D1 _7313_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_15_12 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_15_23 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_85_500 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_15_34 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_85_544 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6709__A2 _6040_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_57_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_38_471 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_53_474 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4520_ _4162_/A _4656_/C _4326_/D _4809_/A vssd2 vssd2 vccd2 vccd2 _4520_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_103_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4451_ _4451_/A _4451_/B vssd2 vssd2 vccd2 vccd2 _4452_/B sky130_fd_sc_hd__xor2_4
Xhold206 wbs_dat_i[3] vssd2 vssd2 vccd2 vccd2 input92/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 _7381_/X vssd2 vssd2 vccd2 vccd2 _7382_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_124 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7170_ _7169_/A _7169_/B _7169_/C vssd2 vssd2 vccd2 vccd2 _7171_/B sky130_fd_sc_hd__a21o_1
Xhold239 _7732_/Q vssd2 vssd2 vccd2 vccd2 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 hold367/X vssd2 vssd2 vccd2 vccd2 _7768_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6121_ _6128_/B _6128_/C vssd2 vssd2 vccd2 vccd2 _6184_/B sky130_fd_sc_hd__nand2_1
XTAP_500 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4382_ _4326_/D _4381_/X _4374_/A _5458_/A vssd2 vssd2 vccd2 vccd2 _4382_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_40_179 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_21_393 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_511 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _6051_/B _6051_/C _6051_/A vssd2 vssd2 vccd2 vccd2 _6052_/Y sky130_fd_sc_hd__a21oi_1
XTAP_544 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5145_/A _5404_/A _4935_/A _4936_/Y _4938_/B vssd2 vssd2 vccd2 vccd2 _5005_/B
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4319__A _4598_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_577 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6954_ _6954_/A _6954_/B vssd2 vssd2 vccd2 vccd2 _6956_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_88_382 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_48_224 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7349__B _7385_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5905_ _5896_/Y _5901_/Y _5903_/Y _5755_/B vssd2 vssd2 vccd2 vccd2 _6783_/A sky130_fd_sc_hd__a31o_4
XFILLER_0_91_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_76_555 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6885_ _6885_/A _6885_/B _6885_/C vssd2 vssd2 vccd2 vccd2 _6887_/A sky130_fd_sc_hd__and3_1
XANTENNA__4054__A _5455_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5836_ _6670_/A _5836_/B _5878_/C vssd2 vssd2 vccd2 vccd2 _5836_/X sky130_fd_sc_hd__and3_1
XFILLER_0_48_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_106_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5767_ _6550_/A vssd2 vssd2 vccd2 vccd2 _5819_/B sky130_fd_sc_hd__inv_2
XFILLER_0_63_249 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4718_ _4718_/A _4718_/B vssd2 vssd2 vccd2 vccd2 _4720_/B sky130_fd_sc_hd__xor2_1
X_7506_ _7565_/A vssd2 vssd2 vccd2 vccd2 _7506_/Y sky130_fd_sc_hd__inv_2
X_5698_ _5694_/A _5694_/B _5694_/C _5694_/D _5735_/B vssd2 vssd2 vccd2 vccd2 _5699_/B
+ sky130_fd_sc_hd__o41a_2
X_4649_ _4649_/A _4649_/B vssd2 vssd2 vccd2 vccd2 _4651_/A sky130_fd_sc_hd__xnor2_2
X_7437_ hold121/X _7799_/D _7451_/S vssd2 vssd2 vccd2 vccd2 _7437_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_97_81 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7368_ _7440_/A _7368_/B vssd2 vssd2 vccd2 vccd2 _7654_/D sky130_fd_sc_hd__and2_1
X_6319_ _6318_/A _6317_/B _7034_/A vssd2 vssd2 vccd2 vccd2 _6393_/A sky130_fd_sc_hd__a21oi_1
X_7299_ _7300_/A _7300_/B vssd2 vssd2 vccd2 vccd2 _7301_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4647__B1 _5406_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_wb_clk_i clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7800_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__6147__C _6705_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_39_213 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_94_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_82_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_94_385 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_82_525 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_67_599 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_109_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_82_569 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_105_384 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_50_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_50_455 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_50_499 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6619__A _7034_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_93_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_26_11 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_58_533 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_58_511 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3951_ _7779_/Q _3954_/C _4050_/B vssd2 vssd2 vccd2 vccd2 _3952_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__6504__D _7237_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_58_566 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_73_536 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6670_ _6670_/A _6670_/B vssd2 vssd2 vccd2 vccd2 _6670_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_45_216 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3882_ _7767_/Q _4326_/B _4144_/D _4267_/D vssd2 vssd2 vccd2 vccd2 _3882_/X sky130_fd_sc_hd__and4_1
XFILLER_0_42_65 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5621_ _5586_/B _5584_/Y _5586_/Y vssd2 vssd2 vccd2 vccd2 _6194_/B sky130_fd_sc_hd__o21a_2
X_5552_ _5530_/B _5532_/B _5530_/A vssd2 vssd2 vccd2 vccd2 _5553_/B sky130_fd_sc_hd__o21bai_1
X_4503_ _4504_/A _4504_/B vssd2 vssd2 vccd2 vccd2 _4558_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_53_293 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5483_ _5483_/A _5483_/B vssd2 vssd2 vccd2 vccd2 _5487_/A sky130_fd_sc_hd__xor2_1
X_4434_ _4863_/A _4704_/B _4711_/A _4782_/B vssd2 vssd2 vccd2 vccd2 _4435_/B sky130_fd_sc_hd__nor4_1
X_7222_ _7222_/A _7222_/B _7222_/C _7294_/C vssd2 vssd2 vccd2 vccd2 _7223_/B sky130_fd_sc_hd__and4_1
X_7153_ _7153_/A _7153_/B vssd2 vssd2 vccd2 vccd2 _7155_/B sky130_fd_sc_hd__xnor2_1
X_4365_ _4348_/A _4348_/B _4346_/Y vssd2 vssd2 vccd2 vccd2 _4372_/A sky130_fd_sc_hd__a21o_1
X_7084_ _7083_/A _7083_/B _7211_/B vssd2 vssd2 vccd2 vccd2 _7131_/C sky130_fd_sc_hd__o21ai_1
X_6104_ _5907_/D _6150_/B _7047_/A _6590_/A vssd2 vssd2 vccd2 vccd2 _6106_/B sky130_fd_sc_hd__a22o_1
XTAP_341 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5152__B _5315_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_385 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _6094_/B _6281_/B _6158_/A _6100_/D vssd2 vssd2 vccd2 vccd2 _6035_/X sky130_fd_sc_hd__and4b_1
X_4296_ _4363_/A _4297_/A vssd2 vssd2 vccd2 vccd2 _4296_/X sky130_fd_sc_hd__and2b_1
XANTENNA__4049__A _7806_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_396 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout283_A _7563_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_95_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_49_500 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1529 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_25 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_36 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_47 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_95_149 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6937_ _6989_/A _7253_/B _6938_/B vssd2 vssd2 vccd2 vccd2 _6937_/X sky130_fd_sc_hd__or3_1
XPHY_58 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_69 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6868_ _6868_/A _6868_/B vssd2 vssd2 vccd2 vccd2 _6869_/B sky130_fd_sc_hd__and2_1
X_5819_ _6436_/A _5819_/B _6402_/A _5907_/D vssd2 vssd2 vccd2 vccd2 _5865_/A sky130_fd_sc_hd__and4_1
XFILLER_0_64_547 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6711__B _7051_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6799_ _6729_/A _6731_/B _6729_/B vssd2 vssd2 vccd2 vccd2 _6808_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_44_271 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_17_496 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_114_181 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_102_321 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_387 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
Xhold581 hold77/X vssd2 vssd2 vccd2 vccd2 input27/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold570 input8/X vssd2 vssd2 vccd2 vccd2 hold86/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 la_data_in[1] vssd2 vssd2 vccd2 vccd2 hold89/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_319 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__3798__A _7768_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_138 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_86_149 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_67_330 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_103_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_55_536 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_82_399 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_50_241 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
Xoutput119 hold643/X vssd2 vssd2 vccd2 vccd2 hold286/A sky130_fd_sc_hd__buf_6
XFILLER_0_105_181 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xoutput108 hold653/X vssd2 vssd2 vccd2 vccd2 hold300/A sky130_fd_sc_hd__buf_6
XANTENNA__6848__A1 _6634_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_11_639 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6349__A _6581_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4150_ _4141_/X _4146_/Y _4147_/Y _4148_/X _3880_/A vssd2 vssd2 vccd2 vccd2 _4155_/A
+ sky130_fd_sc_hd__a41o_1
X_4081_ _4454_/A _4083_/B _4081_/C vssd2 vssd2 vccd2 vccd2 _4081_/X sky130_fd_sc_hd__and3_1
XANTENNA__5823__A2 _7336_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_37_87 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_78_606 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7840_ _7870_/CLK _7840_/D _7599_/Y vssd2 vssd2 vccd2 vccd2 _7840_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_138 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4983_ _4912_/A _4912_/B _4910_/Y vssd2 vssd2 vccd2 vccd2 _4985_/B sky130_fd_sc_hd__a21boi_4
XFILLER_0_58_341 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7771_ _7771_/CLK _7771_/D _7530_/Y vssd2 vssd2 vccd2 vccd2 _7771_/Q sky130_fd_sc_hd__dfrtp_4
X_6722_ _6776_/A _6722_/B vssd2 vssd2 vccd2 vccd2 _6724_/B sky130_fd_sc_hd__and2_1
XANTENNA__6812__A _6812_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3934_ _7783_/Q _3954_/C _3910_/B _4050_/B vssd2 vssd2 vccd2 vccd2 _3935_/B sky130_fd_sc_hd__o31a_2
XFILLER_0_85_193 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6653_ _6582_/A _6582_/C _6582_/B vssd2 vssd2 vccd2 vccd2 _6660_/A sky130_fd_sc_hd__a21boi_2
XFILLER_0_73_322 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_46_558 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3865_ _7761_/Q _4745_/A vssd2 vssd2 vccd2 vccd2 _3865_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_61_517 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5604_ _5612_/B _5606_/C _7866_/Q vssd2 vssd2 vccd2 vccd2 _5828_/B sky130_fd_sc_hd__o21ai_4
X_6584_ _6584_/A _6584_/B vssd2 vssd2 vccd2 vccd2 _6596_/A sky130_fd_sc_hd__nor2_1
X_3796_ _4162_/A vssd2 vssd2 vccd2 vccd2 _4490_/A sky130_fd_sc_hd__inv_2
XANTENNA__4051__B _5455_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5535_ _5535_/A _5535_/B vssd2 vssd2 vccd2 vccd2 _5537_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_641 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_75_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5466_ _5466_/A _5466_/B vssd2 vssd2 vccd2 vccd2 _5470_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7205_ _7205_/A _7205_/B vssd2 vssd2 vccd2 vccd2 _7206_/B sky130_fd_sc_hd__nor2_1
X_4417_ _4417_/A _4417_/B vssd2 vssd2 vccd2 vccd2 _4422_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__3890__B _4162_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5397_ _5398_/A _5398_/B vssd2 vssd2 vccd2 vccd2 _5397_/X sky130_fd_sc_hd__and2b_1
X_7136_ _7104_/A _7104_/B _7102_/Y vssd2 vssd2 vccd2 vccd2 _7155_/A sky130_fd_sc_hd__o21ai_1
X_4348_ _4348_/A _4348_/B vssd2 vssd2 vccd2 vccd2 _4350_/B sky130_fd_sc_hd__xor2_4
X_7067_ _7067_/A _7067_/B vssd2 vssd2 vccd2 vccd2 _7072_/A sky130_fd_sc_hd__xnor2_1
X_4279_ _4221_/A _4220_/A _4220_/B vssd2 vssd2 vccd2 vccd2 _4287_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__4078__A1 _7762_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6018_ _6670_/A _6253_/B _6253_/C _6018_/D vssd2 vssd2 vccd2 vccd2 _6018_/X sky130_fd_sc_hd__and4_1
XFILLER_0_96_447 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_96_425 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1304 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6425__C _6426_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1348 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_119 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4250__A1 _7771_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4250__B2 _4268_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_hold410_A _7886_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_17_293 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_60_583 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_60_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7553__A _7557_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4896__B _5374_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_102_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_87_403 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_90_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_87_469 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_87_447 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6230__A2 _6150_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_300 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_114_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_7_408 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_99_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6351__B _7045_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_43_517 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_113_405 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4152__A _7766_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_70_369 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_3_614 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_113_449 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_23_263 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5320_ _5320_/A _5320_/B vssd2 vssd2 vccd2 vccd2 _5321_/B sky130_fd_sc_hd__nor2_1
X_5251_ _5125_/X _5249_/D _5194_/Y vssd2 vssd2 vccd2 vccd2 _5252_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_48_42 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4202_ _7768_/Q _4519_/B _4519_/C vssd2 vssd2 vccd2 vccd2 _4206_/B sky130_fd_sc_hd__and3_1
X_5182_ _5182_/A _5182_/B vssd2 vssd2 vccd2 vccd2 _5183_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__5414__C _5528_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5133__D _5133_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4133_ _4134_/A _4134_/B vssd2 vssd2 vccd2 vccd2 _4135_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7402__S _7418_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4064_ _7763_/Q _4707_/A _4063_/X _7765_/Q vssd2 vssd2 vccd2 vccd2 _4064_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_64_41 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_64_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7823_ _7826_/CLK _7823_/D _7582_/Y vssd2 vssd2 vccd2 vccd2 _7823_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4046__B _4747_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7638__A _7641_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7754_ _7758_/CLK _7754_/D _7513_/Y vssd2 vssd2 vccd2 vccd2 _7754_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_80_73 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_74_620 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6705_ _6783_/A _6705_/B _7253_/A _7253_/B vssd2 vssd2 vccd2 vccd2 _6706_/B sky130_fd_sc_hd__or4_1
XFILLER_0_58_193 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4966_ _4966_/A _5374_/B vssd2 vssd2 vccd2 vccd2 _4969_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_19_536 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_95 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6509__B1 _7291_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_61_303 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4897_ _4017_/A _4017_/B _5528_/B vssd2 vssd2 vccd2 vccd2 _4899_/B sky130_fd_sc_hd__a21oi_2
X_7685_ _7798_/CLK _7685_/D vssd2 vssd2 vccd2 vccd2 _7685_/Q sky130_fd_sc_hd__dfxtp_1
X_3917_ _7785_/Q _3918_/B vssd2 vssd2 vccd2 vccd2 _4125_/B sky130_fd_sc_hd__xor2_4
X_6636_ _6636_/A _7255_/B vssd2 vssd2 vccd2 vccd2 _6637_/B sky130_fd_sc_hd__nor2_1
X_3848_ _4267_/D _3996_/B vssd2 vssd2 vccd2 vccd2 _4201_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_104_405 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6567_ _6567_/A _6567_/B vssd2 vssd2 vccd2 vccd2 _6604_/A sky130_fd_sc_hd__and2_1
XFILLER_0_89_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5518_ _5518_/A _5518_/B vssd2 vssd2 vccd2 vccd2 _5518_/Y sky130_fd_sc_hd__nand2_1
X_6498_ _6498_/A _6498_/B vssd2 vssd2 vccd2 vccd2 _6500_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__7092__B _7237_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5449_ _5252_/A _5252_/B _5448_/A vssd2 vssd2 vccd2 vccd2 _5449_/Y sky130_fd_sc_hd__a21oi_1
X_7119_ _7072_/A _7072_/B _7066_/X vssd2 vssd2 vccd2 vccd2 _7121_/B sky130_fd_sc_hd__o21a_1
Xfanout187 _6436_/A vssd2 vssd2 vccd2 vccd2 _6590_/A sky130_fd_sc_hd__buf_4
Xfanout198 _4271_/Y vssd2 vssd2 vccd2 vccd2 _5042_/B sky130_fd_sc_hd__clkbuf_8
Xfanout176 _3991_/Y vssd2 vssd2 vccd2 vccd2 _4747_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__6155__C _6253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_96_233 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1112 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_609 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_96_277 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1156 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7548__A _7564_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1189 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_152 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_64_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_25_517 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_25_539 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_100_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_33_572 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6920__B1 _7291_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_110_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_60_391 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_482 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_907 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_288 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_20_299 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_109_69 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA_max_cap211_A _4044_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_18_45 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_18_67 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4462__A1 _4896_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4147__A _7764_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_222 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4462__B2 _4962_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_75_406 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4820_ _4821_/A _4821_/B vssd2 vssd2 vccd2 vccd2 _4820_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_75_439 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__6081__B _6973_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4751_ _4752_/A _4752_/B vssd2 vssd2 vccd2 vccd2 _4751_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_55_152 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_50_32 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_28_344 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_70_111 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4682_ _4683_/B _4683_/A vssd2 vssd2 vccd2 vccd2 _4767_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_50_76 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7470_ _7710_/Q _7483_/A2 _7483_/B1 hold327/X vssd2 vssd2 vccd2 vccd2 _7470_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_28_388 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6421_ _6421_/A _6421_/B vssd2 vssd2 vccd2 vccd2 _6422_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6352_ _6425_/A _6571_/C _6353_/B vssd2 vssd2 vccd2 vccd2 _6352_/X sky130_fd_sc_hd__and3_1
XFILLER_0_59_41 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5303_ _5305_/A _5305_/B vssd2 vssd2 vccd2 vccd2 _5303_/Y sky130_fd_sc_hd__nor2_1
X_6283_ _6283_/A _6283_/B _6587_/B vssd2 vssd2 vccd2 vccd2 _6283_/X sky130_fd_sc_hd__and3_1
XFILLER_0_59_96 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5234_ _5235_/A _5235_/B vssd2 vssd2 vccd2 vccd2 _5295_/B sky130_fd_sc_hd__and2_1
XFILLER_0_11_277 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5165_ _5220_/A _5406_/A vssd2 vssd2 vccd2 vccd2 _5171_/A sky130_fd_sc_hd__or2_1
XFILLER_0_75_73 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA_fanout196_A _4318_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4116_ _4747_/A _5042_/A vssd2 vssd2 vccd2 vccd2 _4118_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_38_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_98_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5096_ _5220_/A _5315_/B vssd2 vssd2 vccd2 vccd2 _5101_/A sky130_fd_sc_hd__nor2_1
X_4047_ _4048_/B vssd2 vssd2 vccd2 vccd2 _4189_/A sky130_fd_sc_hd__inv_2
XPHY_206 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_78_277 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7806_ _7806_/CLK _7806_/D _7565_/Y vssd2 vssd2 vccd2 vccd2 _7806_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__7368__A _7440_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_38_108 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XPHY_228 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5998_ _5998_/A _5998_/B _5998_/C vssd2 vssd2 vccd2 vccd2 _6001_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_47_620 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4205__B2 _7767_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4205__A1 _7765_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_81_409 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4949_ _4949_/A _4949_/B _4949_/C vssd2 vssd2 vccd2 vccd2 _4950_/B sky130_fd_sc_hd__nor3_1
X_7737_ _7739_/CLK _7737_/D _7496_/Y vssd2 vssd2 vccd2 vccd2 _7737_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_366 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7668_ _7779_/CLK _7668_/D vssd2 vssd2 vccd2 vccd2 _7668_/Q sky130_fd_sc_hd__dfxtp_1
X_6619_ _7034_/A _6769_/B vssd2 vssd2 vccd2 vccd2 _6620_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_61_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4508__A2 _5222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_34_347 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7599_ _7627_/A vssd2 vssd2 vccd2 vccd2 _7599_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_69_211 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_97_586 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_97_597 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_38_675 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_37_152 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_111_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_20_24 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_20_46 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_21_542 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XTAP_704 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_66 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_726 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6970_ _6970_/A _7033_/D vssd2 vssd2 vccd2 vccd2 _7826_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_45_43 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5921_ _6074_/A _6071_/B _6019_/C _5921_/D vssd2 vssd2 vccd2 vccd2 _5923_/C sky130_fd_sc_hd__and4_1
XANTENNA__6092__A _6092_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_75_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_75_214 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5852_ _6253_/A _6100_/D _6587_/B _5938_/C vssd2 vssd2 vccd2 vccd2 _5853_/C sky130_fd_sc_hd__and4_1
X_4803_ _4803_/A _4803_/B _4803_/C vssd2 vssd2 vccd2 vccd2 _4804_/B sky130_fd_sc_hd__and3_1
XFILLER_0_61_75 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5783_ _6093_/A _5850_/B _5936_/B _5850_/D vssd2 vssd2 vccd2 vccd2 _5783_/X sky130_fd_sc_hd__and4_1
XFILLER_0_28_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4734_ _4088_/A _4088_/B _5374_/B vssd2 vssd2 vccd2 vccd2 _4737_/A sky130_fd_sc_hd__a21oi_1
X_7522_ _7524_/A vssd2 vssd2 vccd2 vccd2 _7522_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7137__B1 _7222_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_44_645 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_114_533 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_71_464 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4665_ _4017_/A _4017_/B _5374_/B vssd2 vssd2 vccd2 vccd2 _4668_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_43_155 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7453_ _7350_/C _7453_/B _7453_/C vssd2 vssd2 vccd2 vccd2 _7453_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_0_16_369 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6404_ _6707_/A _6634_/B _6404_/C _6404_/D vssd2 vssd2 vccd2 vccd2 _6405_/B sky130_fd_sc_hd__and4b_1
XANTENNA_fanout209_A _4807_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7384_ _7450_/A _7384_/B vssd2 vssd2 vccd2 vccd2 _7662_/D sky130_fd_sc_hd__and2_1
XFILLER_0_12_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4596_ _4594_/X _4595_/X _4252_/B vssd2 vssd2 vccd2 vccd2 _5326_/B sky130_fd_sc_hd__o21a_1
X_6335_ _6335_/A _6335_/B vssd2 vssd2 vccd2 vccd2 _6337_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_101_205 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_101_81 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_101_249 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6266_ _6855_/A _6973_/A vssd2 vssd2 vccd2 vccd2 _6267_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_86_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6197_ _6550_/A _6479_/C vssd2 vssd2 vccd2 vccd2 _6199_/C sky130_fd_sc_hd__nor2_1
X_5217_ _5217_/A _5217_/B vssd2 vssd2 vccd2 vccd2 _5219_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__5871__B1 _7846_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5148_ _4250_/X _4251_/X _4256_/X _5030_/C _4214_/C vssd2 vssd2 vccd2 vccd2 _5149_/B
+ sky130_fd_sc_hd__o311a_1
XANTENNA__6415__A2 _6989_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5079_ _5079_/A _5079_/B vssd2 vssd2 vccd2 vccd2 _5089_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4426__A1 _4162_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4426__B2 _7772_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_109_305 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_66_236 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5926__A1 _7844_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_109_349 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6730__A _7037_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_34_100 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__5926__B2 _7845_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_62_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_22_306 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_34_177 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6639__C1 _5992_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6654__A2 _7094_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5081__A _5210_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_89_317 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_106_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6811__C1 _7294_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5614__B1 _5645_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_350 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_15_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_85_523 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_57_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_85_556 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_72_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_25_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_26_645 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_38_494 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_53_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5256__A _5548_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_41_615 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4450_ _4451_/A _4451_/B vssd2 vssd2 vccd2 vccd2 _4450_/Y sky130_fd_sc_hd__nor2_1
Xhold207 input92/X vssd2 vssd2 vccd2 vccd2 hold207/X sky130_fd_sc_hd__buf_1
XFILLER_0_25_188 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
Xwire171 _5860_/Y vssd2 vssd2 vccd2 vccd2 _6138_/A sky130_fd_sc_hd__clkbuf_4
Xhold229 _7737_/Q vssd2 vssd2 vccd2 vccd2 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 hold375/X vssd2 vssd2 vccd2 vccd2 _7762_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4381_ _7772_/Q _4458_/D _4326_/B _4809_/A vssd2 vssd2 vccd2 vccd2 _4381_/X sky130_fd_sc_hd__a22o_1
X_6120_ _6119_/B _6119_/C _6119_/A vssd2 vssd2 vccd2 vccd2 _6128_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_383 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_501 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6087__A _6707_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6051_ _6051_/A _6051_/B _6051_/C vssd2 vssd2 vccd2 vccd2 _6051_/X sky130_fd_sc_hd__and3_1
XTAP_545 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _4951_/A _4951_/B _4950_/A vssd2 vssd2 vccd2 vccd2 _5005_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_42 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_578 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7410__S _7418_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6953_ _6954_/A _6954_/B vssd2 vssd2 vccd2 vccd2 _7010_/B sky130_fd_sc_hd__and2_1
XFILLER_0_72_85 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6884_ _6919_/B _6883_/C _6883_/A vssd2 vssd2 vccd2 vccd2 _6885_/C sky130_fd_sc_hd__a21o_1
X_5904_ _5896_/Y _5901_/Y _5903_/Y _5755_/B vssd2 vssd2 vccd2 vccd2 _6634_/B sky130_fd_sc_hd__a31oi_4
X_5835_ _6253_/B _6253_/C _6018_/D _5835_/D vssd2 vssd2 vccd2 vccd2 _5878_/C sky130_fd_sc_hd__and4_1
XFILLER_0_76_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_8_355 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_8_344 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_29_461 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_29_483 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_91_548 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6550__A _6550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_44_431 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5766_ hold415/X _5761_/X _5765_/Y _5845_/B vssd2 vssd2 vccd2 vccd2 _6550_/A sky130_fd_sc_hd__o2bb2a_4
X_4717_ _4717_/A _4717_/B vssd2 vssd2 vccd2 vccd2 _4718_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_44_464 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7505_ _7565_/A vssd2 vssd2 vccd2 vccd2 _7505_/Y sky130_fd_sc_hd__inv_2
X_5697_ _7884_/Q _5697_/B vssd2 vssd2 vccd2 vccd2 _6100_/D sky130_fd_sc_hd__xnor2_4
XANTENNA__4173__C_N _5030_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_102_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_71_272 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4648_ _4649_/A _4649_/B vssd2 vssd2 vccd2 vccd2 _4648_/Y sky130_fd_sc_hd__nand2_1
X_7436_ _7436_/A _7436_/B vssd2 vssd2 vccd2 vccd2 _7686_/D sky130_fd_sc_hd__and2_1
XFILLER_0_16_188 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4070__A _4328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_31_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4579_ _4580_/A _4580_/B vssd2 vssd2 vccd2 vccd2 _4579_/Y sky130_fd_sc_hd__nand2_1
X_7367_ hold139/X _7766_/D _7383_/S vssd2 vssd2 vccd2 vccd2 _7367_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6318_ _6318_/A _6318_/B vssd2 vssd2 vccd2 vccd2 _7817_/D sky130_fd_sc_hd__xnor2_1
X_7298_ _7316_/A _7298_/B vssd2 vssd2 vccd2 vccd2 _7300_/B sky130_fd_sc_hd__and2b_1
XANTENNA__6097__B1 _6670_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6249_ _6311_/C _6249_/B vssd2 vssd2 vccd2 vccd2 _6316_/B sky130_fd_sc_hd__xor2_1
XANTENNA__6147__D _6939_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_79_350 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_39_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_109_113 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6163__C _7094_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7556__A _7557_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5076__A _5145_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_22_147 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7291__A _7291_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_22_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_101_591 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__6088__B1 _5948_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_26_23 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_89_125 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold90 hold90/A vssd2 vssd2 vccd2 vccd2 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_169 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_58_523 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_3950_ _7778_/Q _3950_/B vssd2 vssd2 vccd2 vccd2 _4018_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_42_11 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_58_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_58_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3881_ _7765_/Q _3886_/C _4144_/C vssd2 vssd2 vccd2 vccd2 _3881_/X sky130_fd_sc_hd__and3_1
XFILLER_0_73_548 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_45_239 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5620_ _7846_/Q _5620_/B _5620_/C _6075_/C vssd2 vssd2 vccd2 vccd2 _5620_/X sky130_fd_sc_hd__and4_1
XFILLER_0_53_250 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5551_ _4809_/B _4814_/Y _5529_/B _5550_/Y vssd2 vssd2 vccd2 vccd2 _5553_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_81_570 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4502_ _4502_/A _4502_/B vssd2 vssd2 vccd2 vccd2 _4504_/B sky130_fd_sc_hd__xnor2_2
X_7221_ _7291_/A _7253_/B _7253_/C _7253_/A vssd2 vssd2 vccd2 vccd2 _7223_/A sky130_fd_sc_hd__o22a_1
X_5482_ _5483_/A _5483_/B vssd2 vssd2 vccd2 vccd2 _5515_/B sky130_fd_sc_hd__nand2b_1
X_4433_ _5042_/A _4711_/A _4782_/B _4863_/A vssd2 vssd2 vccd2 vccd2 _4433_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_0_67_30 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7152_ _7152_/A _7152_/B vssd2 vssd2 vccd2 vccd2 _7153_/B sky130_fd_sc_hd__xor2_1
X_4364_ _4356_/A _4356_/B _4354_/Y vssd2 vssd2 vccd2 vccd2 _4415_/A sky130_fd_sc_hd__a21oi_2
X_7083_ _7083_/A _7083_/B _7211_/B vssd2 vssd2 vccd2 vccd2 _7131_/B sky130_fd_sc_hd__or3_1
XFILLER_0_67_52 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_342 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6103_ _6093_/X _6098_/X _6101_/X _6102_/X _5769_/B vssd2 vssd2 vccd2 vccd2 _6103_/X
+ sky130_fd_sc_hd__o41a_2
X_4295_ _4236_/X _4239_/B _4235_/X vssd2 vssd2 vccd2 vccd2 _4363_/A sky130_fd_sc_hd__a21oi_2
XTAP_375 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ _6282_/A _5937_/B _5938_/C _6094_/B _6157_/A vssd2 vssd2 vccd2 vccd2 _6034_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_386 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6545__A _6707_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_83_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA_fanout276_A _7454_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_20_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_68_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1508 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1519 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6936_ _7047_/A _7222_/A vssd2 vssd2 vccd2 vccd2 _6938_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_49_523 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_15 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_26 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_37 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_49_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_9_620 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XPHY_48 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_59 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_76_386 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6867_ _6868_/A _6868_/B vssd2 vssd2 vccd2 vccd2 _6916_/A sky130_fd_sc_hd__nor2_1
XANTENNA__7376__A _7452_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5818_ _5868_/B vssd2 vssd2 vccd2 vccd2 _5818_/Y sky130_fd_sc_hd__inv_2
X_6798_ _6798_/A _6798_/B vssd2 vssd2 vccd2 vccd2 _6826_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_559 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_36_228 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_91_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5749_ _3803_/Y _6094_/B _6510_/B _6283_/B vssd2 vssd2 vccd2 vccd2 _5749_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_0_72_570 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_44_283 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_32_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_114_193 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_102_333 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7419_ _7452_/A _7419_/B vssd2 vssd2 vccd2 vccd2 _7678_/D sky130_fd_sc_hd__and2_1
XFILLER_0_4_380 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold571 hold86/X vssd2 vssd2 vccd2 vccd2 _7855_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold560 la_data_in[28] vssd2 vssd2 vccd2 vccd2 hold73/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_399 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold582 input27/X vssd2 vssd2 vccd2 vccd2 hold78/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 hold89/X vssd2 vssd2 vccd2 vccd2 input12/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5997__C _6855_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5045__A1 _5220_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_82_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_55_515 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_103_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6190__A _7336_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_82_345 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__7337__A3 _6669_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_12_36 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_113_609 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_70_529 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_88_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_23_467 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_105_193 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xoutput109 hold671/X vssd2 vssd2 vccd2 vccd2 hold318/A sky130_fd_sc_hd__buf_6
XANTENNA__6848__A2 _7197_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6349__B _6989_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_37_22 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4080_ _4519_/C _4267_/C _4201_/D _4080_/D vssd2 vssd2 vccd2 vccd2 _4081_/C sky130_fd_sc_hd__and4_1
X_4982_ _4982_/A _4982_/B vssd2 vssd2 vccd2 vccd2 _4985_/A sky130_fd_sc_hd__xnor2_4
X_7770_ _7787_/CLK _7770_/D _7529_/Y vssd2 vssd2 vccd2 vccd2 _7770_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_92_109 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7814_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_6721_ _6721_/A _6721_/B vssd2 vssd2 vccd2 vccd2 _6722_/B sky130_fd_sc_hd__or2_1
XANTENNA__6812__B _6812_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_46_504 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3933_ _3954_/C _3910_/B _4050_/B vssd2 vssd2 vccd2 vccd2 _3936_/B sky130_fd_sc_hd__o21ai_2
X_6652_ _6572_/D _6652_/B vssd2 vssd2 vccd2 vccd2 _6661_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_73_334 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_46_537 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_46_548 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_3864_ _4082_/B _4201_/D _3864_/C vssd2 vssd2 vccd2 vccd2 _3864_/X sky130_fd_sc_hd__and3_1
XFILLER_0_33_209 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5603_ _5612_/B _5606_/C _7866_/Q vssd2 vssd2 vccd2 vccd2 _5607_/A sky130_fd_sc_hd__o21a_1
X_6583_ _6582_/A _6582_/B _6582_/C vssd2 vssd2 vccd2 vccd2 _6584_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_14_412 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3795_ _7771_/Q vssd2 vssd2 vccd2 vccd2 _4521_/A sky130_fd_sc_hd__inv_2
X_5534_ _5535_/B _5535_/A vssd2 vssd2 vccd2 vccd2 _5534_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_41_220 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5971__A1_N _7336_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_78_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5465_ _5465_/A _5465_/B vssd2 vssd2 vccd2 vccd2 _5466_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7204_ _7205_/A _7205_/B vssd2 vssd2 vccd2 vccd2 _7246_/B sky130_fd_sc_hd__and2_1
XFILLER_0_68_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4416_ _4417_/A _4417_/B vssd2 vssd2 vccd2 vccd2 _4480_/A sky130_fd_sc_hd__nand2_1
X_7135_ _7326_/A _7326_/B _7034_/A vssd2 vssd2 vccd2 vccd2 _7174_/A sky130_fd_sc_hd__a21oi_1
X_5396_ _5398_/B _5398_/A vssd2 vssd2 vccd2 vccd2 _5396_/Y sky130_fd_sc_hd__nand2b_1
X_4347_ _4347_/A _4347_/B vssd2 vssd2 vccd2 vccd2 _4348_/B sky130_fd_sc_hd__xor2_4
X_7066_ _7067_/A _7067_/B vssd2 vssd2 vccd2 vccd2 _7066_/X sky130_fd_sc_hd__or2_1
XANTENNA__4078__A2 _4809_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4278_ _4882_/A _4896_/A _4226_/A _4227_/Y vssd2 vssd2 vccd2 vccd2 _4289_/A sky130_fd_sc_hd__o31ai_4
XFILLER_0_94_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6275__A _6812_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6017_ _6157_/A _6017_/B vssd2 vssd2 vccd2 vccd2 _6017_/X sky130_fd_sc_hd__and2_1
XTAP_1305 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_128 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6224__B1 _6152_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_96_459 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1338 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_364 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6919_ _6919_/A _6919_/B vssd2 vssd2 vccd2 vccd2 _6928_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_52_529 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_17_261 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_60_573 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_141 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_32_297 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold390 _7655_/Q vssd2 vssd2 vccd2 vccd2 hold390/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4710__B1 _5099_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_415 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_59_128 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_114_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_28_515 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5140__A2_N _5431_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_23_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_83_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_99_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_36_570 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_113_417 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_82_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_11_404 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_23_242 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5250_ _5250_/A _5250_/B _5250_/C _5250_/D vssd2 vssd2 vccd2 vccd2 _5252_/A sky130_fd_sc_hd__or4_1
XFILLER_0_23_286 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__5264__A _5315_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4201_ _4809_/A _4519_/C _4267_/C _4201_/D vssd2 vssd2 vccd2 vccd2 _4206_/A sky130_fd_sc_hd__and4_1
X_5181_ _5182_/A _5182_/B vssd2 vssd2 vccd2 vccd2 _5181_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_54 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5414__D _5528_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4132_ _4132_/A _4132_/B vssd2 vssd2 vccd2 vccd2 _4134_/B sky130_fd_sc_hd__xnor2_1
X_4063_ _4252_/D _4063_/B _4252_/B vssd2 vssd2 vccd2 vccd2 _4063_/X sky130_fd_sc_hd__and3b_1
X_7822_ _7826_/CLK _7822_/D _7581_/Y vssd2 vssd2 vccd2 vccd2 _7822_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4046__C _4898_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_673 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4965_ _5220_/A _4965_/B vssd2 vssd2 vccd2 vccd2 _4970_/A sky130_fd_sc_hd__or2_2
X_7753_ _7758_/CLK _7753_/D _7512_/Y vssd2 vssd2 vccd2 vccd2 _7753_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_63 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6704_ _6705_/B _7253_/A _7253_/B _6783_/A vssd2 vssd2 vccd2 vccd2 _6704_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6509__A1 _5816_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3916_ _7786_/Q _3916_/B vssd2 vssd2 vccd2 vccd2 _4252_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_19_548 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4896_ _4896_/A _5374_/B vssd2 vssd2 vccd2 vccd2 _4899_/A sky130_fd_sc_hd__or2_2
X_7684_ _7800_/CLK _7684_/D vssd2 vssd2 vccd2 vccd2 _7684_/Q sky130_fd_sc_hd__dfxtp_1
X_6635_ _6635_/A _6635_/B vssd2 vssd2 vccd2 vccd2 _6637_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_73_186 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7182__A1 _7181_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3847_ _7797_/Q _3847_/B vssd2 vssd2 vccd2 vccd2 _4148_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_417 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6566_ _6566_/A _6566_/B _6566_/C vssd2 vssd2 vccd2 vccd2 _6567_/B sky130_fd_sc_hd__or3_1
XFILLER_0_61_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__4997__B _4997_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_6_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_14_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5517_ _5517_/A vssd2 vssd2 vccd2 vccd2 _5561_/A sky130_fd_sc_hd__inv_2
X_6497_ _6939_/A _6572_/B vssd2 vssd2 vccd2 vccd2 _6498_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_14_275 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5448_ _5448_/A vssd2 vssd2 vccd2 vccd2 _5448_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7485__A2 _7453_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5379_ _5379_/A _5379_/B vssd2 vssd2 vccd2 vccd2 _5380_/B sky130_fd_sc_hd__nor2_1
X_7118_ _7166_/B _7120_/B vssd2 vssd2 vccd2 vccd2 _7121_/A sky130_fd_sc_hd__nor2_1
XANTENNA__5902__A _6093_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xfanout188 _5674_/X vssd2 vssd2 vccd2 vccd2 _6436_/A sky130_fd_sc_hd__buf_2
Xfanout199 _4271_/Y vssd2 vssd2 vccd2 vccd2 _5145_/A sky130_fd_sc_hd__clkbuf_4
Xfanout177 _4708_/A vssd2 vssd2 vccd2 vccd2 _4598_/A sky130_fd_sc_hd__buf_6
X_7049_ _6357_/X _6359_/X _6281_/B _7143_/B vssd2 vssd2 vccd2 vccd2 _7052_/A sky130_fd_sc_hd__o211a_1
XANTENNA__6436__C _7222_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4518__A _4736_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_96_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XTAP_1113 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_437 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_96_289 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_84_407 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1146 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4253__A _7768_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_64_131 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_52_304 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_37_378 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_64_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_52_359 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7564__A _7564_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_18_592 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_33_551 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_20_201 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_103_494 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XTAP_908 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7476__A2 _7483_/A2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_20_267 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_919 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5812__A _6093_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4147__B _4809_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_34_56 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_34_78 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6362__B _7099_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_68_481 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4750_ _4601_/A _4601_/B _4669_/B _4670_/B _4670_/A vssd2 vssd2 vccd2 vccd2 _4752_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_11 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_28_356 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4163__A _4268_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_83_473 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_71_613 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4681_ _4681_/A _4681_/B vssd2 vssd2 vccd2 vccd2 _4683_/B sky130_fd_sc_hd__xor2_1
X_6420_ _6421_/A _6421_/B vssd2 vssd2 vccd2 vccd2 _6420_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_70_123 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_50_88 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_113_225 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6351_ _6812_/A _7045_/A vssd2 vssd2 vccd2 vccd2 _6353_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5706__B _6670_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5302_ _5139_/A _5139_/B _5243_/B _5242_/B _5242_/A vssd2 vssd2 vccd2 vccd2 _5305_/B
+ sky130_fd_sc_hd__a32oi_4
XANTENNA__7467__A2 _7454_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6282_ _6282_/A _6510_/B vssd2 vssd2 vccd2 vccd2 _6282_/X sky130_fd_sc_hd__and2_1
X_5233_ _5233_/A _5233_/B vssd2 vssd2 vccd2 vccd2 _5235_/B sky130_fd_sc_hd__xor2_1
X_5164_ _5164_/A _5164_/B vssd2 vssd2 vccd2 vccd2 _5176_/A sky130_fd_sc_hd__nor2_1
XANTENNA__5722__A _6152_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4115_ _4104_/X _4108_/X _4115_/C _4115_/D vssd2 vssd2 vccd2 vccd2 _4704_/B sky130_fd_sc_hd__and4bb_4
X_5095_ _5160_/A _5095_/B vssd2 vssd2 vccd2 vccd2 _5111_/A sky130_fd_sc_hd__nor2_2
XANTENNA_fanout189_A _5142_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4046_ _4598_/A _4747_/A _4898_/A _4882_/A vssd2 vssd2 vccd2 vccd2 _4048_/B sky130_fd_sc_hd__or4_1
XFILLER_0_91_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_78_245 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XPHY_207 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7805_ _7806_/CLK _7805_/D _7564_/Y vssd2 vssd2 vccd2 vccd2 _7805_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_229 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_218 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_93_237 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5997_ _6105_/A _6105_/B _6855_/A _6939_/A vssd2 vssd2 vccd2 vccd2 _5998_/C sky130_fd_sc_hd__or4_1
X_4948_ _4949_/A _4949_/B _4949_/C vssd2 vssd2 vccd2 vccd2 _4950_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_74_451 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_46_131 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_46_120 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7736_ _7739_/CLK _7736_/D _7495_/Y vssd2 vssd2 vccd2 vccd2 _7736_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4073__A _7765_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4879_ _4810_/A _4811_/A _5498_/D _4808_/A _4808_/B vssd2 vssd2 vccd2 vccd2 _4887_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_62_613 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_101 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_46_153 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7667_ _7779_/CLK _7667_/D vssd2 vssd2 vccd2 vccd2 _7667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_315 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_34_326 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6618_ _6467_/B _6618_/B vssd2 vssd2 vccd2 vccd2 _6769_/B sky130_fd_sc_hd__and2b_1
XANTENNA__5166__B1 _4814_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_46_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7384__A _7450_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_34_359 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_15_540 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7598_ _7627_/A vssd2 vssd2 vccd2 vccd2 _7598_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5931__A_N _6550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6549_ _6670_/A _7313_/A vssd2 vssd2 vccd2 vccd2 _6549_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_42_381 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_30_521 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7458__A2 _7454_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6728__A _6973_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_100_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7091__B1 _7222_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7559__A _7563_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_84_226 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_57_429 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_65_440 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_37_164 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_111_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_108_586 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_443 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__4711__A _4711_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_52_134 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_25_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5807__A _6253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_80_498 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_21_521 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_96_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_705 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_45_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5920_ _6398_/A _5921_/D _5979_/D _5920_/D vssd2 vssd2 vccd2 vccd2 _5923_/B sky130_fd_sc_hd__and4_1
XFILLER_0_48_418 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6092__B _6939_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_61_43 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5851_ _7845_/Q _6281_/B _5700_/Y _6283_/B _7843_/Q vssd2 vssd2 vccd2 vccd2 _5851_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_259 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4802_ _4803_/A _4803_/B _4803_/C vssd2 vssd2 vccd2 vccd2 _4804_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__4199__B2 _4162_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4199__A1 _4656_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5782_ _6282_/A _5936_/B _5936_/C vssd2 vssd2 vccd2 vccd2 _5782_/X sky130_fd_sc_hd__and3_1
XANTENNA__7137__A1 _7099_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4733_ _4733_/A _4733_/B vssd2 vssd2 vccd2 vccd2 _4753_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_304 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7521_ _7557_/A vssd2 vssd2 vccd2 vccd2 _7521_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_164 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_29_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_114_501 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7137__B2 _6430_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_56_495 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_43_123 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7408__S _7418_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7452_ _7452_/A _7452_/B vssd2 vssd2 vccd2 vccd2 _7694_/D sky130_fd_sc_hd__and2_1
XFILLER_0_28_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_114_545 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6403_ _6783_/A _6479_/C _7051_/A _6707_/A vssd2 vssd2 vccd2 vccd2 _6405_/A sky130_fd_sc_hd__o22a_1
X_4664_ _4664_/A _4664_/B vssd2 vssd2 vccd2 vccd2 _4670_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_668 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_71_487 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7383_ hold146/X _7662_/Q _7383_/S vssd2 vssd2 vccd2 vccd2 _7383_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_510 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_381 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__3882__D _4267_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4595_ _4809_/A _4030_/B _4427_/A _7771_/Q _4815_/B vssd2 vssd2 vccd2 vccd2 _4595_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_114_589 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6334_ _6335_/A _6334_/B vssd2 vssd2 vccd2 vccd2 _6412_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_101_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6265_ _6634_/B _6571_/B vssd2 vssd2 vccd2 vccd2 _6267_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6548__A _6670_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5216_ _5216_/A _5216_/B vssd2 vssd2 vccd2 vccd2 _5217_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_50_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4123__A1 _4328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6196_ _7143_/A vssd2 vssd2 vccd2 vccd2 _6479_/C sky130_fd_sc_hd__inv_2
XANTENNA__5871__A1 _6670_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4068__A _7762_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5147_ _4314_/X _4317_/X _4954_/C _4214_/B vssd2 vssd2 vccd2 vccd2 _5149_/A sky130_fd_sc_hd__o211a_1
XFILLER_0_98_307 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5078_ _5168_/A _5145_/B vssd2 vssd2 vccd2 vccd2 _5079_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_79_543 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4029_ _4315_/B _4427_/A _4164_/C _4036_/B vssd2 vssd2 vccd2 vccd2 _4029_/X sky130_fd_sc_hd__and4_1
XANTENNA__6283__A _6283_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_79_565 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_79_554 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_39_429 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_109_317 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_81_207 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7719_ _7750_/CLK _7719_/D vssd2 vssd2 vccd2 vccd2 _7719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_501 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_62_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6730__B _7045_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_62_454 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6639__B1 _7143_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5362__A _5404_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5081__B _5210_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5311__B1 _5550_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_89_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_106_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6811__B1 _6664_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_57_215 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_72_229 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_53_410 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_31_46 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_80_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_31_79 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_53_487 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6878__B1 _7222_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold208 _7394_/X vssd2 vssd2 vccd2 vccd2 _7395_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_178 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_40_104 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold219 _7359_/X vssd2 vssd2 vccd2 vccd2 _7360_/B sky130_fd_sc_hd__dlygate4sd3_1
X_4380_ _4454_/A _4380_/B vssd2 vssd2 vccd2 vccd2 _4380_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_40_159 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_111_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_502 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6087__B _6581_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6050_ _6049_/A _6049_/B _6049_/C vssd2 vssd2 vccd2 vccd2 _6051_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_56_21 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XTAP_535 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _5128_/A _4996_/B _4992_/Y vssd2 vssd2 vccd2 vccd2 _5068_/A sky130_fd_sc_hd__a21o_1
XTAP_568 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_98 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4319__C _4782_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_88_362 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_76_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6952_ _6952_/A _6952_/B vssd2 vssd2 vccd2 vccd2 _6954_/B sky130_fd_sc_hd__xnor2_1
X_6883_ _6883_/A _6919_/B _6883_/C vssd2 vssd2 vccd2 vccd2 _6885_/B sky130_fd_sc_hd__nand3_1
X_5903_ _6282_/A _5769_/X _5785_/X _6157_/A _5902_/X vssd2 vssd2 vccd2 vccd2 _5903_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_72_97 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5834_ _6019_/D _5834_/B _5834_/C vssd2 vssd2 vccd2 vccd2 _5834_/X sky130_fd_sc_hd__and3_1
XFILLER_0_91_527 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_91_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_106_309 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6550__B _7255_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_56_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5765_ _5992_/C _5853_/A _5762_/X _5764_/X vssd2 vssd2 vccd2 vccd2 _5765_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_0_16_112 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_98_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4716_ _4717_/A _4717_/B vssd2 vssd2 vccd2 vccd2 _4716_/X sky130_fd_sc_hd__or2_1
XFILLER_0_71_240 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA_fanout221_A _5081_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7504_ _7565_/A vssd2 vssd2 vccd2 vccd2 _7504_/Y sky130_fd_sc_hd__inv_2
X_5696_ _7884_/Q _5697_/B vssd2 vssd2 vccd2 vccd2 _6283_/B sky130_fd_sc_hd__xor2_4
X_4647_ wire212/X _4881_/A2 _5406_/A vssd2 vssd2 vccd2 vccd2 _4649_/B sky130_fd_sc_hd__a21oi_2
X_7435_ hold139/X _7686_/Q _7451_/S vssd2 vssd2 vccd2 vccd2 _7435_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_126 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7366_ _7436_/A _7366_/B vssd2 vssd2 vccd2 vccd2 _7653_/D sky130_fd_sc_hd__and2_1
X_6317_ _7034_/A _6317_/B vssd2 vssd2 vccd2 vccd2 _6318_/B sky130_fd_sc_hd__nor2_1
X_4578_ wire212/X _4881_/A2 _5315_/B vssd2 vssd2 vccd2 vccd2 _4580_/B sky130_fd_sc_hd__a21oi_2
X_7297_ _7297_/A _7297_/B _7297_/C vssd2 vssd2 vccd2 vccd2 _7298_/B sky130_fd_sc_hd__or3_1
XANTENNA__6097__A1 _7847_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6248_ _6186_/A _6186_/B _6184_/X vssd2 vssd2 vccd2 vccd2 _6249_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__6097__B2 _7846_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6179_ _6180_/B _6180_/A vssd2 vssd2 vccd2 vccd2 _6308_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__4526__A _4810_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_94_321 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_67_557 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_39_248 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_109_125 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_109_169 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_35_432 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_35_454 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__5076__B _5328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7572__A _7613_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4335__A1 _4863_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_22_137 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7291__B _7291_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6088__A1 _6634_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7285__B1 _7336_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6088__B2 _5931_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5820__A _7886_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_89_137 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold91 hold91/A vssd2 vssd2 vccd2 vccd2 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 hold80/A vssd2 vssd2 vccd2 vccd2 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_181 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_58_557 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6155__A_N _6152_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_85_387 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_73_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_45_207 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3880_ _3880_/A _4002_/B _4002_/C _3880_/D vssd2 vssd2 vccd2 vccd2 _3880_/X sky130_fd_sc_hd__and4_1
XFILLER_0_45_229 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_26_421 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5550_ _5550_/A _5550_/B vssd2 vssd2 vccd2 vccd2 _5550_/Y sky130_fd_sc_hd__nor2_1
X_4501_ _4502_/A _4502_/B vssd2 vssd2 vccd2 vccd2 _4501_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_13_104 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5481_ _5515_/A _5481_/B vssd2 vssd2 vccd2 vccd2 _5483_/B sky130_fd_sc_hd__and2_1
X_7220_ _7310_/A _7220_/B vssd2 vssd2 vccd2 vccd2 _7831_/D sky130_fd_sc_hd__xnor2_1
X_4432_ _5042_/A _4711_/A _4782_/B _4863_/A vssd2 vssd2 vccd2 vccd2 _4435_/A sky130_fd_sc_hd__o22a_1
XFILLER_0_41_446 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_41_457 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7151_ _7152_/A _7152_/B vssd2 vssd2 vccd2 vccd2 _7151_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1_576 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4363_ _4363_/A _4418_/B _4297_/A vssd2 vssd2 vccd2 vccd2 _4417_/A sky130_fd_sc_hd__nor3b_2
X_7082_ _7082_/A _7082_/B vssd2 vssd2 vccd2 vccd2 _7211_/B sky130_fd_sc_hd__or2_1
XTAP_321 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6102_ _6253_/A _6102_/B _6102_/C vssd2 vssd2 vccd2 vccd2 _6102_/X sky130_fd_sc_hd__and3_1
X_4294_ _4294_/A _4294_/B vssd2 vssd2 vccd2 vccd2 _4297_/A sky130_fd_sc_hd__xor2_2
X_6033_ _6092_/A _6855_/A vssd2 vssd2 vccd2 vccd2 _6045_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_67_97 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_376 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7421__S _7451_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6545__B _7253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_107_81 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1509 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6935_ _6039_/X _6040_/X _7222_/C _5992_/B vssd2 vssd2 vccd2 vccd2 _6938_/A sky130_fd_sc_hd__o211a_1
XFILLER_0_49_513 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XPHY_16 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_38 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_76_321 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XPHY_49 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_76_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_76_354 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_64_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6866_ _6866_/A _6866_/B vssd2 vssd2 vccd2 vccd2 _6868_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5817_ _6436_/A _6402_/A _5907_/D _5819_/B vssd2 vssd2 vccd2 vccd2 _5868_/B sky130_fd_sc_hd__a22o_1
X_6797_ _6797_/A _6797_/B vssd2 vssd2 vccd2 vccd2 _6798_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_91_368 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4081__A _4454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_17_465 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5748_ _7843_/Q _6281_/B _5747_/Y _7844_/Q _6094_/B vssd2 vssd2 vccd2 vccd2 _5748_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_72_582 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_17_476 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5679_ _5694_/A _5694_/B _5694_/C _5735_/B vssd2 vssd2 vccd2 vccd2 _5679_/X sky130_fd_sc_hd__o31a_1
XANTENNA__4317__A1 _4268_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_102_345 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7418_ hold146/X _7790_/D _7418_/S vssd2 vssd2 vccd2 vccd2 _7418_/X sky130_fd_sc_hd__mux2_1
X_7349_ _7349_/A _7385_/B vssd2 vssd2 vccd2 vccd2 _7349_/Y sky130_fd_sc_hd__nand2_1
Xhold572 la_data_in[4] vssd2 vssd2 vccd2 vccd2 hold79/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold550 input15/X vssd2 vssd2 vccd2 vccd2 hold72/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 hold73/X vssd2 vssd2 vccd2 vccd2 input21/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 hold78/X vssd2 vssd2 vccd2 vccd2 _7840_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 input12/X vssd2 vssd2 vccd2 vccd2 hold90/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5817__B2 _5819_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_99_424 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__5997__D _6939_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5045__A2 _4965_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7567__A _7613_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_67_321 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_12_59 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_12_48 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_112_109 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_105_161 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5815__A _5816_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_23_435 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_23_457 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_50_287 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5550__A _5550_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_77_118 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_98_490 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4981_ _4981_/A _4981_/B vssd2 vssd2 vccd2 vccd2 _4982_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_58_321 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_85_162 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6720_ _6721_/A _6721_/B vssd2 vssd2 vccd2 vccd2 _6776_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6812__C _7253_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_58_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_46_516 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3932_ _4252_/B _4125_/B _4252_/D _4707_/A vssd2 vssd2 vccd2 vccd2 _4315_/B sky130_fd_sc_hd__nor4_4
X_6651_ _6651_/A _6651_/B vssd2 vssd2 vccd2 vccd2 _6685_/A sky130_fd_sc_hd__and2_1
X_3863_ _4268_/A _4083_/B _3901_/B vssd2 vssd2 vccd2 vccd2 _3864_/C sky130_fd_sc_hd__and3_1
X_6582_ _6582_/A _6582_/B _6582_/C vssd2 vssd2 vccd2 vccd2 _6584_/A sky130_fd_sc_hd__and3_1
XFILLER_0_73_368 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5602_ _5645_/B _7865_/Q vssd2 vssd2 vccd2 vccd2 _5606_/C sky130_fd_sc_hd__and2_2
XFILLER_0_54_582 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_6_668 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5533_ _5500_/A _5500_/B _5463_/A vssd2 vssd2 vccd2 vccd2 _5535_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__6941__C1 _6152_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3794_ _4268_/A vssd2 vssd2 vccd2 vccd2 _4457_/A sky130_fd_sc_hd__inv_2
XFILLER_0_81_390 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5725__A _6152_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7416__S _7418_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_41_210 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_112_621 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_14_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5464_ _5465_/A _5465_/B vssd2 vssd2 vccd2 vccd2 _5466_/A sky130_fd_sc_hd__or2_1
XFILLER_0_112_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_78_85 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7203_ _7203_/A _7203_/B vssd2 vssd2 vccd2 vccd2 _7205_/B sky130_fd_sc_hd__xor2_1
X_5395_ _5395_/A _5395_/B vssd2 vssd2 vccd2 vccd2 _5398_/B sky130_fd_sc_hd__nand2_2
X_4415_ _4415_/A _4415_/B vssd2 vssd2 vccd2 vccd2 _4417_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_41_287 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7134_ _7134_/A _7134_/B vssd2 vssd2 vccd2 vccd2 _7326_/B sky130_fd_sc_hd__nor2_1
X_4346_ _4347_/A _4347_/B vssd2 vssd2 vccd2 vccd2 _4346_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6556__A _6556_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7065_ _7005_/A _7005_/B _6981_/X vssd2 vssd2 vccd2 vccd2 _7067_/B sky130_fd_sc_hd__a21oi_1
X_4277_ _4277_/A _4277_/B vssd2 vssd2 vccd2 vccd2 _4291_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__6275__B _6812_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6472__B2 _6670_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3899__B _7768_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6016_ _7849_/Q _6016_/B _6071_/B vssd2 vssd2 vccd2 vccd2 _6016_/X sky130_fd_sc_hd__and3_1
XFILLER_0_68_118 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1339 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_490 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1317 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_376 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6918_ _6738_/A _7313_/B _6669_/X _6664_/A vssd2 vssd2 vccd2 vccd2 _6930_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_37_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6849_ _6795_/A _6795_/B _6792_/Y vssd2 vssd2 vccd2 vccd2 _6871_/A sky130_fd_sc_hd__a21o_1
XANTENNA__5906__A2_N _6707_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_17_240 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_32_210 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_32_232 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_103_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_102_153 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_20_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_32_287 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4710__A1 _5042_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold380 _7652_/Q vssd2 vssd2 vccd2 vccd2 hold380/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4710__B2 _4711_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold391 hold692/X vssd2 vssd2 vccd2 vccd2 _7786_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_67_151 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_23_14 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_23_25 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_67_195 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_23_47 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_28_549 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_82_121 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_55_346 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_113_429 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_51_530 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7479__B1 _7483_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_11_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5264__B _5374_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4200_ _4268_/A _4200_/B vssd2 vssd2 vccd2 vccd2 _4200_/X sky130_fd_sc_hd__and2_1
X_5180_ _5111_/A _5111_/B _5109_/X vssd2 vssd2 vccd2 vccd2 _5182_/B sky130_fd_sc_hd__a21oi_2
X_4131_ _4132_/A _4132_/B vssd2 vssd2 vccd2 vccd2 _4181_/A sky130_fd_sc_hd__and2b_1
X_4062_ _4060_/Y _4061_/X _4707_/A vssd2 vssd2 vccd2 vccd2 _4062_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_427 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_78_416 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7821_ _7826_/CLK _7821_/D _7580_/Y vssd2 vssd2 vccd2 vccd2 _7821_/Q sky130_fd_sc_hd__dfrtp_1
X_4964_ _5033_/A _4964_/B vssd2 vssd2 vccd2 vccd2 _4974_/A sky130_fd_sc_hd__and2_2
X_7752_ _7758_/CLK _7752_/D _7511_/Y vssd2 vssd2 vccd2 vccd2 _7752_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4046__D _4882_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6703_ _6661_/A _6661_/B _6659_/X vssd2 vssd2 vccd2 vccd2 _6721_/A sky130_fd_sc_hd__a21o_1
X_3915_ _7785_/Q _3954_/C _3910_/B _3907_/X _4050_/B vssd2 vssd2 vccd2 vccd2 _3916_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_0_19_516 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_19_527 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6509__A2 _5816_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4895_ _5099_/A _5220_/A vssd2 vssd2 vccd2 vccd2 _4900_/A sky130_fd_sc_hd__nor2_2
X_7683_ _7795_/CLK _7683_/D vssd2 vssd2 vccd2 vccd2 _7683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_508 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6634_ _6707_/A _6634_/B _7222_/A _7222_/C vssd2 vssd2 vccd2 vccd2 _6635_/B sky130_fd_sc_hd__and4b_1
XFILLER_0_73_176 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7182__A2 _7253_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3846_ _7797_/Q _3847_/B vssd2 vssd2 vccd2 vccd2 _3996_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_27_582 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6565_ _6566_/A _6566_/B _6566_/C vssd2 vssd2 vccd2 vccd2 _6567_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_80_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_54_390 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_42_541 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_42_530 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6496_ _6496_/A _6496_/B vssd2 vssd2 vccd2 vccd2 _6498_/A sky130_fd_sc_hd__xor2_1
XANTENNA__5455__A _5455_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5516_ _5516_/A _5516_/B vssd2 vssd2 vccd2 vccd2 _5517_/A sky130_fd_sc_hd__nor2_1
X_5447_ _5447_/A _5447_/B _5445_/A _5445_/B vssd2 vssd2 vccd2 vccd2 _5448_/A sky130_fd_sc_hd__or4bb_2
XFILLER_0_42_585 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7092__D _7253_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5454__C_N _5547_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5378_ _5381_/A vssd2 vssd2 vccd2 vccd2 _5412_/B sky130_fd_sc_hd__inv_2
X_7117_ _7117_/A _7117_/B vssd2 vssd2 vccd2 vccd2 _7120_/B sky130_fd_sc_hd__nor2_1
X_4329_ _7767_/Q _4656_/C _4893_/B _7766_/Q vssd2 vssd2 vccd2 vccd2 _4329_/X sky130_fd_sc_hd__a22o_1
Xfanout167 _6082_/A vssd2 vssd2 vccd2 vccd2 _6402_/A sky130_fd_sc_hd__buf_4
X_7048_ _7048_/A _7048_/B vssd2 vssd2 vccd2 vccd2 _7058_/A sky130_fd_sc_hd__xor2_1
Xfanout178 _7138_/C vssd2 vssd2 vccd2 vccd2 _7253_/A sky130_fd_sc_hd__buf_4
Xfanout189 _5142_/C vssd2 vssd2 vccd2 vccd2 _5404_/A sky130_fd_sc_hd__buf_4
XANTENNA__4518__B _5220_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_416 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1114 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1147 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd2 vssd2 vccd2 vccd2 clkbuf_leaf_9_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_482 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1169 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_184 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_37_324 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_37_346 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_37_357 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_107_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_64_176 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_52_316 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_18_560 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_80_658 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_100_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4931__A1 _4779_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_909 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_27 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6196__A _7143_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_18_25 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5812__B _6424_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_87_202 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_87_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_56_611 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_55_110 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4680_ _4681_/B _4681_/A vssd2 vssd2 vccd2 vccd2 _4680_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_519 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_71_669 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_70_135 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_113_237 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6350_ _6664_/A _7047_/A vssd2 vssd2 vccd2 vccd2 _6353_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_168 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_24_541 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5301_ _5301_/A _5301_/B vssd2 vssd2 vccd2 vccd2 _5305_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_213 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__3919__C_N _7764_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_76 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6281_ _6510_/A _6281_/B _6281_/C vssd2 vssd2 vccd2 vccd2 _6281_/X sky130_fd_sc_hd__and3_2
XFILLER_0_59_87 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5232_ _5233_/A _5233_/B vssd2 vssd2 vccd2 vccd2 _5295_/A sky130_fd_sc_hd__and2_1
X_5163_ _5163_/A _5163_/B vssd2 vssd2 vccd2 vccd2 _5183_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_53 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4114_ _4109_/X _4112_/X _4113_/X _4103_/A vssd2 vssd2 vccd2 vccd2 _4115_/C sky130_fd_sc_hd__a31o_1
X_5094_ _4172_/Y _5164_/B _5550_/B _4129_/Y vssd2 vssd2 vccd2 vccd2 _5095_/B sky130_fd_sc_hd__o22a_1
X_4045_ _4747_/A _4898_/A _4882_/A _4598_/A vssd2 vssd2 vccd2 vccd2 _4053_/B sky130_fd_sc_hd__o22ai_1
XFILLER_0_78_213 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_93_205 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA_fanout251_A _6069_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7804_ _7804_/CLK _7804_/D _7563_/Y vssd2 vssd2 vccd2 vccd2 _7804_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_219 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_208 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5996_ _5907_/D _5948_/X _5994_/X _6590_/A vssd2 vssd2 vccd2 vccd2 _5998_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_19_313 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_93_249 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4947_ _4947_/A _4947_/B vssd2 vssd2 vccd2 vccd2 _4949_/C sky130_fd_sc_hd__xor2_1
X_7735_ _7739_/CLK _7735_/D _7494_/Y vssd2 vssd2 vccd2 vccd2 _7735_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_463 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4878_ _4801_/A _4801_/B _4798_/X vssd2 vssd2 vccd2 vccd2 _4889_/A sky130_fd_sc_hd__a21bo_1
X_7666_ _7779_/CLK _7666_/D vssd2 vssd2 vccd2 vccd2 _7666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_305 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6617_ _6765_/A _6617_/B vssd2 vssd2 vccd2 vccd2 _6769_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_187 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_3829_ _4745_/A _4454_/B _4656_/C _4006_/B vssd2 vssd2 vccd2 vccd2 _4458_/C sky130_fd_sc_hd__or4_4
X_7597_ _7597_/A vssd2 vssd2 vccd2 vccd2 _7597_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_552 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_61_179 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6548_ _6670_/A _7313_/A vssd2 vssd2 vccd2 vccd2 _7294_/B sky130_fd_sc_hd__and2_1
XFILLER_0_30_500 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6479_ _6783_/A _6855_/A _6479_/C _7051_/A vssd2 vssd2 vccd2 vccd2 _6481_/B sky130_fd_sc_hd__or4_1
XFILLER_0_30_544 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_30_577 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6728__B _6973_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7091__A1 _6430_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7091__B2 _7197_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_268 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_65_463 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_20_15 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_111_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_80_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4711__B _5042_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_53_669 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_21_555 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_103_281 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_706 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_79 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_88_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_45_67 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5850_ _6510_/A _5850_/B _5936_/B _5850_/D vssd2 vssd2 vccd2 vccd2 _5857_/A sky130_fd_sc_hd__and4_1
X_4801_ _4801_/A _4801_/B vssd2 vssd2 vccd2 vccd2 _4803_/C sky130_fd_sc_hd__xnor2_1
X_5781_ _6670_/B _5781_/B _6358_/B vssd2 vssd2 vccd2 vccd2 _5936_/C sky130_fd_sc_hd__and3b_1
X_4732_ _4732_/A _4732_/B vssd2 vssd2 vccd2 vccd2 _4733_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_56_452 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7520_ _7557_/A vssd2 vssd2 vccd2 vccd2 _7520_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7137__A2 _7222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4663_ _4663_/A _4663_/B vssd2 vssd2 vccd2 vccd2 _4664_/B sky130_fd_sc_hd__nand2_1
X_7451_ hold146/X _7806_/D _7451_/S vssd2 vssd2 vccd2 vccd2 _7451_/X sky130_fd_sc_hd__mux2_1
X_6402_ _6402_/A _7145_/A vssd2 vssd2 vccd2 vccd2 _6406_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_71_499 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7382_ _7452_/A _7382_/B vssd2 vssd2 vccd2 vccd2 _7661_/D sky130_fd_sc_hd__and2_1
X_4594_ _7772_/Q _4019_/Y _4032_/C _4656_/A vssd2 vssd2 vccd2 vccd2 _4594_/X sky130_fd_sc_hd__a22o_1
X_6333_ _6335_/B vssd2 vssd2 vccd2 vccd2 _6334_/B sky130_fd_sc_hd__inv_2
XFILLER_0_12_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_12_544 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6264_ _6217_/A _6216_/A _6216_/B vssd2 vssd2 vccd2 vccd2 _6271_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_86_41 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5215_ _5216_/A _5216_/B vssd2 vssd2 vccd2 vccd2 _5215_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_86_85 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6195_ _6191_/X _6192_/X _6193_/X _6194_/X _5630_/B vssd2 vssd2 vccd2 vccd2 _6404_/C
+ sky130_fd_sc_hd__o41a_4
X_5146_ _5146_/A _5146_/B vssd2 vssd2 vccd2 vccd2 _5158_/A sky130_fd_sc_hd__xnor2_1
X_5077_ _5077_/A _5077_/B vssd2 vssd2 vccd2 vccd2 _5079_/A sky130_fd_sc_hd__nand2_1
X_4028_ _4706_/A1 _3965_/A _3986_/X _7767_/Q _4162_/B vssd2 vssd2 vccd2 vccd2 _4028_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_109_329 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5979_ _6670_/A _6194_/B _6019_/D _5979_/D vssd2 vssd2 vccd2 vccd2 _5979_/X sky130_fd_sc_hd__and4_1
XFILLER_0_19_110 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4812__A _5042_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7718_ _7750_/CLK _7718_/D vssd2 vssd2 vccd2 vccd2 _7718_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__7395__A _7440_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_19_165 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_62_411 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7649_ _7795_/CLK _7649_/D vssd2 vssd2 vccd2 vccd2 _7649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_488 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_15_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6639__A1 _6039_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_100_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6404__A_N _6707_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5362__B _5406_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5311__A1 _5276_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5311__B2 _5210_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5081__C _5081_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5075__B1 _5076_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_15_48 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_65_260 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_31_25 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_108_395 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_53_466 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6878__A1 _6571_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6878__B2 _6571_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_111_505 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold209 hold383/X vssd2 vssd2 vccd2 vccd2 _7793_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_503 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5133_/A _5133_/B _5548_/A vssd2 vssd2 vccd2 vccd2 _5069_/A sky130_fd_sc_hd__a21oi_1
XTAP_536 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7055__A1 _7140_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3801__A _6093_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6951_ _6952_/A _6952_/B vssd2 vssd2 vccd2 vccd2 _7010_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_76_525 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5902_ _6093_/A _5936_/B _5936_/C vssd2 vssd2 vccd2 vccd2 _5902_/X sky130_fd_sc_hd__and3_1
X_6882_ _6881_/A _6919_/A _6881_/C vssd2 vssd2 vccd2 vccd2 _6883_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_76_569 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_76_547 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_29_430 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5833_ _6398_/A _6071_/B _6424_/A vssd2 vssd2 vccd2 vccd2 _5834_/C sky130_fd_sc_hd__and3_1
XANTENNA__4632__A _4704_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_8_324 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_17_614 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_44_400 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_7503_ _7565_/A vssd2 vssd2 vccd2 vccd2 _7503_/Y sky130_fd_sc_hd__inv_2
X_5764_ _6102_/B _6102_/C _5764_/C vssd2 vssd2 vccd2 vccd2 _5764_/X sky130_fd_sc_hd__and3_1
XFILLER_0_29_496 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4715_ _4636_/A _4633_/X _4635_/B vssd2 vssd2 vccd2 vccd2 _4717_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_71_252 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_44_444 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5695_ _7883_/Q _5694_/X _5735_/B vssd2 vssd2 vccd2 vccd2 _5697_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_114_321 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_71_285 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4646_ _5029_/A _5222_/A vssd2 vssd2 vccd2 vccd2 _4649_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_44_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7434_ _7436_/A _7434_/B vssd2 vssd2 vccd2 vccd2 _7685_/D sky130_fd_sc_hd__and2_1
XANTENNA_fanout214_A _6404_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_31_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_114_365 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_102_527 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_102_516 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_71_296 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4577_ _5029_/A _4965_/B vssd2 vssd2 vccd2 vccd2 _4580_/A sky130_fd_sc_hd__nor2_1
X_7365_ hold169/X _7765_/D _7383_/S vssd2 vssd2 vccd2 vccd2 _7365_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_102_538 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_97_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6316_ _6316_/A _6316_/B vssd2 vssd2 vccd2 vccd2 _6317_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_12_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7296_ _7297_/A _7297_/B _7297_/C vssd2 vssd2 vccd2 vccd2 _7316_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_110_593 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6247_ _6308_/B _6247_/B vssd2 vssd2 vccd2 vccd2 _6311_/C sky130_fd_sc_hd__xnor2_2
X_6178_ _6119_/A _6119_/C _6119_/B vssd2 vssd2 vccd2 vccd2 _6180_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_99_617 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5129_ _4996_/B _5249_/C _5250_/C _5250_/A vssd2 vssd2 vccd2 vccd2 _5130_/B sky130_fd_sc_hd__o2bb2a_2
XANTENNA__4807__A _4807_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4526__B _5315_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_67_503 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_94_333 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_109_137 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_82_517 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5638__A _6158_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_94_399 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_75_580 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5357__B _5357_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_90_550 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_62_241 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_47_293 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_35_466 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5076__C _5404_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_62_274 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_50_425 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_7_390 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_50_447 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_15_190 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_30_160 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_30_171 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6088__A2 _6664_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6493__C1 _5992_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_89_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
Xhold70 hold70/A vssd2 vssd2 vccd2 vccd2 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 hold81/A vssd2 vssd2 vccd2 vccd2 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A vssd2 vssd2 vccd2 vccd2 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_149 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_97_193 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_85_322 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_73_517 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5548__A _5548_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5771__A1 _6283_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_26_433 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_81_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4500_ _4500_/A _4500_/B vssd2 vssd2 vccd2 vccd2 _4502_/B sky130_fd_sc_hd__xor2_2
X_5480_ _5480_/A _5480_/B _5480_/C vssd2 vssd2 vccd2 vccd2 _5481_/B sky130_fd_sc_hd__or3_1
XFILLER_0_101_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4431_ _4598_/A _5276_/A vssd2 vssd2 vccd2 vccd2 _4436_/A sky130_fd_sc_hd__nor2_2
XANTENNA_1 _7385_/Y vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_111_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5283__A _5431_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7150_ _7152_/A _7152_/B vssd2 vssd2 vccd2 vccd2 _7191_/B sky130_fd_sc_hd__and2_1
X_4362_ _4362_/A _4362_/B vssd2 vssd2 vccd2 vccd2 _7734_/D sky130_fd_sc_hd__xnor2_1
X_7081_ _7081_/A _7081_/B _7081_/C vssd2 vssd2 vccd2 vccd2 _7082_/B sky130_fd_sc_hd__nor3_2
XTAP_322 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6101_ _6099_/X _6100_/X _5850_/B vssd2 vssd2 vccd2 vccd2 _6101_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_21_193 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4293_ _4293_/A _4293_/B vssd2 vssd2 vccd2 vccd2 _4294_/B sky130_fd_sc_hd__xnor2_2
X_6032_ _6032_/A _6032_/B vssd2 vssd2 vccd2 vccd2 _6051_/A sky130_fd_sc_hd__xor2_1
XTAP_366 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5039__B1 _5550_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_107_93 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6934_ _6885_/A _6885_/C _6885_/B vssd2 vssd2 vccd2 vccd2 _6952_/A sky130_fd_sc_hd__a21boi_1
XPHY_17 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_28 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_39 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5458__A _5458_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6865_ _6865_/A _6865_/B vssd2 vssd2 vccd2 vccd2 _6866_/B sky130_fd_sc_hd__xor2_1
X_5816_ _5816_/A _5816_/B vssd2 vssd2 vccd2 vccd2 _5907_/D sky130_fd_sc_hd__nand2_4
X_6796_ _6797_/B _6797_/A vssd2 vssd2 vccd2 vccd2 _6796_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_57_580 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_36_219 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5747_ _5691_/A _5691_/B _6155_/B vssd2 vssd2 vccd2 vccd2 _5747_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_44_263 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_32_403 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5678_ _7877_/Q _7878_/Q vssd2 vssd2 vccd2 vccd2 _5694_/C sky130_fd_sc_hd__or2_2
X_7417_ _7450_/A _7417_/B vssd2 vssd2 vccd2 vccd2 _7677_/D sky130_fd_sc_hd__and2_1
X_4629_ _4708_/A _4736_/A _5142_/C _5076_/D vssd2 vssd2 vccd2 vccd2 _4699_/A sky130_fd_sc_hd__or4_2
XFILLER_0_102_357 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_7348_ _7453_/B _7436_/A _7385_/B hold99/X vssd2 vssd2 vccd2 vccd2 _7348_/X sky130_fd_sc_hd__and4_1
Xhold551 hold72/X vssd2 vssd2 vccd2 vccd2 _7861_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 input21/X vssd2 vssd2 vccd2 vccd2 hold74/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold540 la_data_in[29] vssd2 vssd2 vccd2 vccd2 hold63/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_379 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7279_ _7279_/A _7279_/B vssd2 vssd2 vccd2 vccd2 _7279_/Y sky130_fd_sc_hd__nand2_1
Xhold584 la_data_in[7] vssd2 vssd2 vccd2 vccd2 hold83/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 hold79/X vssd2 vssd2 vccd2 vccd2 input43/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 hold90/X vssd2 vssd2 vccd2 vccd2 _7872_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5817__A2 _6402_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_99_447 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_67_344 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_94_141 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_67_377 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4272__A _4810_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_82_369 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_35_230 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5815__B _5816_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_23_425 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_23_447 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_50_299 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__5550__B _5550_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6662__A _6664_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4980_ _4981_/A _4981_/B vssd2 vssd2 vccd2 vccd2 _4980_/X sky130_fd_sc_hd__and2b_1
X_3931_ _4252_/B _4252_/D vssd2 vssd2 vccd2 vccd2 _3931_/Y sky130_fd_sc_hd__nor2_1
X_6650_ _6650_/A _6650_/B vssd2 vssd2 vccd2 vccd2 _6651_/B sky130_fd_sc_hd__or2_1
XFILLER_0_58_388 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_3862_ _3858_/A _3858_/B _4100_/B _3993_/D vssd2 vssd2 vccd2 vccd2 _3901_/B sky130_fd_sc_hd__a211oi_2
X_6581_ _6581_/A _7140_/A vssd2 vssd2 vccd2 vccd2 _6582_/C sky130_fd_sc_hd__nor2_1
X_5601_ _5581_/A _5581_/B _5581_/C _5579_/X _5645_/B vssd2 vssd2 vccd2 vccd2 _5612_/B
+ sky130_fd_sc_hd__o41a_4
XFILLER_0_54_572 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_5_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5532_ _5532_/A _5532_/B vssd2 vssd2 vccd2 vccd2 _5535_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_263 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6941__B1 _7143_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3793_ _4656_/A vssd2 vssd2 vccd2 vccd2 _3893_/B sky130_fd_sc_hd__inv_2
XFILLER_0_14_436 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_26_296 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5463_ _5463_/A _5463_/B _5526_/A vssd2 vssd2 vccd2 vccd2 _5465_/B sky130_fd_sc_hd__or3b_1
X_7202_ _7203_/A _7203_/B vssd2 vssd2 vccd2 vccd2 _7246_/A sky130_fd_sc_hd__nor2_1
X_5394_ _5394_/A _5394_/B vssd2 vssd2 vccd2 vccd2 _5398_/A sky130_fd_sc_hd__xnor2_4
X_4414_ _4415_/A _4415_/B vssd2 vssd2 vccd2 vccd2 _4479_/A sky130_fd_sc_hd__or2_1
XFILLER_0_41_299 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7133_ _7134_/A _7133_/B vssd2 vssd2 vccd2 vccd2 _7829_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_97 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4345_ _4345_/A _4345_/B vssd2 vssd2 vccd2 vccd2 _4347_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_10_675 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_94_41 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7064_ _7064_/A _7064_/B vssd2 vssd2 vccd2 vccd2 _7067_/A sky130_fd_sc_hd__xnor2_1
X_4276_ _4276_/A _4276_/B vssd2 vssd2 vccd2 vccd2 _4277_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_94_85 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6275__C _6989_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6015_ _7846_/Q _7313_/A _6398_/B _7847_/Q vssd2 vssd2 vccd2 vccd2 _6015_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4483__A1 _5455_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_fanout281_A _7557_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6572__A _6989_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1329 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd2 vssd2 vccd2 vccd2 clkbuf_leaf_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6917_ _7019_/A _6916_/X _6855_/A _7291_/B vssd2 vssd2 vccd2 vccd2 _6961_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_91_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6848_ _6634_/B _7197_/B _6964_/A _6847_/X vssd2 vssd2 vccd2 vccd2 _6897_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_49_399 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_49_388 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_9_430 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_64_347 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_52_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_107_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6779_ _6734_/A _6734_/B _6732_/X vssd2 vssd2 vccd2 vccd2 _6797_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_32_266 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_102_121 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_13_480 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_32_277 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_102_165 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold370 _7670_/Q vssd2 vssd2 vccd2 vccd2 hold370/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 _7667_/Q vssd2 vssd2 vccd2 vccd2 hold381/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4710__A2 _4782_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold392 hold691/X vssd2 vssd2 vccd2 vccd2 _7789_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4267__A _4656_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_28_506 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_43_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_wb_clk_i clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7771_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_328 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5826__A _6158_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_36_550 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_63_391 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_23_222 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_51_553 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_23_233 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6151__A1 _5816_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_2_149 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__6657__A _7047_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4130_ _4598_/A _5029_/A vssd2 vssd2 vccd2 vccd2 _4132_/B sky130_fd_sc_hd__nor2_1
X_4061_ _4252_/B _4252_/C _4252_/D _7766_/Q vssd2 vssd2 vccd2 vccd2 _4061_/X sky130_fd_sc_hd__or4b_1
XANTENNA__4280__C_N _5030_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7820_ _7826_/CLK _7820_/D _7579_/Y vssd2 vssd2 vccd2 vccd2 _7820_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_450 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4963_ _5164_/A _5406_/A _5164_/B _4962_/A vssd2 vssd2 vccd2 vccd2 _4964_/B sky130_fd_sc_hd__o22ai_1
X_7751_ _7758_/CLK _7751_/D _7510_/Y vssd2 vssd2 vccd2 vccd2 _7751_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_54 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6702_ _6645_/A _6645_/B _6646_/X vssd2 vssd2 vccd2 vccd2 _6724_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_58_185 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_3914_ _3954_/C _3910_/B _3907_/X _7790_/Q vssd2 vssd2 vccd2 vccd2 _3918_/B sky130_fd_sc_hd__o31a_2
X_7682_ _7795_/CLK _7682_/D vssd2 vssd2 vccd2 vccd2 _7682_/Q sky130_fd_sc_hd__dfxtp_1
X_6633_ _6783_/A _7253_/A _7253_/B _6707_/A vssd2 vssd2 vccd2 vccd2 _6635_/A sky130_fd_sc_hd__o22a_1
XFILLER_0_74_645 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4894_ _4810_/A _5550_/B _4958_/A _4891_/Y vssd2 vssd2 vccd2 vccd2 _4904_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_46_336 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5717__A1 _6157_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_104_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7427__S _7451_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3845_ _4267_/D vssd2 vssd2 vccd2 vccd2 _4141_/D sky130_fd_sc_hd__inv_2
X_6564_ _6564_/A _6564_/B vssd2 vssd2 vccd2 vccd2 _6566_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_61_328 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_6_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6495_ _6989_/A _6973_/B _6496_/B vssd2 vssd2 vccd2 vccd2 _6495_/X sky130_fd_sc_hd__or3_1
XFILLER_0_42_553 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5515_ _5515_/A _5515_/B _5515_/C vssd2 vssd2 vccd2 vccd2 _5516_/B sky130_fd_sc_hd__and3_1
XFILLER_0_73_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5446_ _5352_/X _5396_/Y _5445_/X _5354_/X _5397_/X vssd2 vssd2 vccd2 vccd2 _5451_/A
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_100_658 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_10_472 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5377_ _5377_/A _5377_/B vssd2 vssd2 vccd2 vccd2 _5381_/A sky130_fd_sc_hd__xnor2_2
X_7116_ _7117_/A _7117_/B vssd2 vssd2 vccd2 vccd2 _7166_/B sky130_fd_sc_hd__and2_1
X_4328_ _4328_/A _4328_/B vssd2 vssd2 vccd2 vccd2 _4328_/X sky130_fd_sc_hd__and2_1
Xfanout168 _6215_/C vssd2 vssd2 vccd2 vccd2 _6939_/A sky130_fd_sc_hd__buf_4
X_7047_ _7047_/A _7294_/B vssd2 vssd2 vccd2 vccd2 _7048_/B sky130_fd_sc_hd__nand2_1
Xfanout179 _6642_/B vssd2 vssd2 vccd2 vccd2 _7181_/A sky130_fd_sc_hd__buf_6
X_4259_ _4260_/A _4260_/B _4260_/C vssd2 vssd2 vccd2 vccd2 _4356_/A sky130_fd_sc_hd__o21a_1
XTAP_1104 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_428 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4815__A _4893_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1137 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_461 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1159 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_271 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_18_550 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_25_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_107_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_64_188 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_52_328 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4931__A2 _5431_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_60_361 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_109_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_18_48 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_87_225 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_87_214 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__4725__A _5029_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4444__B _4966_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_83_420 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_56_645 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_28_325 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_43_317 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_113_205 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_113_249 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5300_ _5300_/A _5300_/B vssd2 vssd2 vccd2 vccd2 _5301_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_51_361 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6280_ _5816_/A _5816_/B _7140_/A vssd2 vssd2 vccd2 vccd2 _6289_/A sky130_fd_sc_hd__a21oi_2
X_5231_ _5231_/A _5231_/B vssd2 vssd2 vccd2 vccd2 _5233_/B sky130_fd_sc_hd__xor2_1
X_5162_ _5162_/A _5162_/B _5162_/C vssd2 vssd2 vccd2 vccd2 _5163_/B sky130_fd_sc_hd__nand3_1
X_5093_ _5093_/A _5093_/B vssd2 vssd2 vccd2 vccd2 _5115_/A sky130_fd_sc_hd__xor2_4
X_4113_ _4374_/A _4149_/B _4149_/C vssd2 vssd2 vccd2 vccd2 _4113_/X sky130_fd_sc_hd__or3_1
XFILLER_0_75_65 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4044_ _4044_/A _4044_/B vssd2 vssd2 vccd2 vccd2 _4882_/A sky130_fd_sc_hd__and2_4
XFILLER_0_78_269 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7803_ _7806_/CLK _7803_/D _7562_/Y vssd2 vssd2 vccd2 vccd2 _7803_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_209 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_93_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5995_ _5991_/X _5993_/X _5781_/B vssd2 vssd2 vccd2 vccd2 _6215_/C sky130_fd_sc_hd__o21ai_2
X_7734_ _7739_/CLK _7734_/D _7493_/Y vssd2 vssd2 vccd2 vccd2 _7734_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3949__B1 _4050_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4946_ _4946_/A _4946_/B vssd2 vssd2 vccd2 vccd2 _4947_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4877_ _4877_/A _4877_/B vssd2 vssd2 vccd2 vccd2 _4912_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_46_166 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7665_ _7779_/CLK _7665_/D vssd2 vssd2 vccd2 vccd2 _7665_/Q sky130_fd_sc_hd__dfxtp_1
X_7596_ _7597_/A vssd2 vssd2 vccd2 vccd2 _7596_/Y sky130_fd_sc_hd__inv_2
X_6616_ _6462_/B _6615_/Y _6765_/B vssd2 vssd2 vccd2 vccd2 _6617_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_15_520 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3828_ _4745_/A _4454_/B _4656_/C _4893_/B vssd2 vssd2 vccd2 vccd2 _4519_/C sky130_fd_sc_hd__nor4_4
X_6547_ _6547_/A _6547_/B vssd2 vssd2 vccd2 vccd2 _6551_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_61_147 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_6_274 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_15_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_391 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6478_ _5948_/X _6404_/C _6404_/D _6634_/B vssd2 vssd2 vccd2 vccd2 _6481_/A sky130_fd_sc_hd__a22o_1
X_5429_ _5430_/A _5430_/B vssd2 vssd2 vccd2 vccd2 _5483_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_100_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6728__C _7140_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5626__B1 _5645_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4429__A1 _4328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7091__A2 _7222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_69_236 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_69_225 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_97_567 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_108_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_65_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_80_412 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7294__C _7294_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_37_199 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4711__C _4782_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_52_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_40_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_80_489 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_21_501 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_33_350 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_293 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_707 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_88_556 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_88_589 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4800_ _5030_/A _5030_/B _4800_/C vssd2 vssd2 vccd2 vccd2 _4801_/B sky130_fd_sc_hd__and3_1
XANTENNA__6042__B1 _5992_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_wire212_A _4044_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6593__A1 _6668_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6670__A _6670_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5780_ _6281_/B _6281_/C vssd2 vssd2 vccd2 vccd2 _5780_/X sky130_fd_sc_hd__and2_1
XTAP_1490 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_209 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4731_ _4732_/A _4732_/B vssd2 vssd2 vccd2 vccd2 _4731_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_56_464 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4662_ _4807_/A _4662_/B _5099_/A _5315_/B vssd2 vssd2 vccd2 vccd2 _4663_/B sky130_fd_sc_hd__or4_1
X_7450_ _7450_/A _7450_/B vssd2 vssd2 vccd2 vccd2 _7693_/D sky130_fd_sc_hd__and2_1
X_6401_ _6550_/A _7253_/A vssd2 vssd2 vccd2 vccd2 _6410_/A sky130_fd_sc_hd__or2_2
XFILLER_0_101_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4593_ _4593_/A _4593_/B vssd2 vssd2 vccd2 vccd2 _4603_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7381_ hold212/X _7773_/D _7383_/S vssd2 vssd2 vccd2 vccd2 _7381_/X sky130_fd_sc_hd__mux2_1
X_6332_ _6332_/A _6332_/B vssd2 vssd2 vccd2 vccd2 _6335_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_523 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6263_ _6138_/A _6973_/B _6206_/B _6207_/X vssd2 vssd2 vccd2 vccd2 _6272_/A sky130_fd_sc_hd__o31ai_4
XFILLER_0_86_53 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5214_ _5149_/A _5149_/B _5153_/A vssd2 vssd2 vccd2 vccd2 _5216_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_86_97 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6194_ _6253_/A _6194_/B _6194_/C vssd2 vssd2 vccd2 vccd2 _6194_/X sky130_fd_sc_hd__and3_1
X_5145_ _5145_/A _5145_/B _5146_/A vssd2 vssd2 vccd2 vccd2 _5201_/B sky130_fd_sc_hd__or3_2
XFILLER_0_36_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_98_309 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5076_ _5145_/A _5328_/A _5404_/A _5076_/D vssd2 vssd2 vccd2 vccd2 _5077_/B sky130_fd_sc_hd__or4_1
X_4027_ _4814_/B _4063_/B _5030_/A vssd2 vssd2 vccd2 vccd2 _4066_/D sky130_fd_sc_hd__and3_1
XFILLER_0_94_526 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_66_228 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_94_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6580__A _6812_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5978_ _6282_/A _6194_/C _6130_/C vssd2 vssd2 vccd2 vccd2 _5978_/X sky130_fd_sc_hd__and3_1
X_4929_ _4930_/A _4930_/B vssd2 vssd2 vccd2 vccd2 _5064_/A sky130_fd_sc_hd__nor2_2
XANTENNA__4812__B _5220_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7717_ _7750_/CLK _7717_/D vssd2 vssd2 vccd2 vccd2 _7717_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4595__B1 _7771_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7648_ _7793_/CLK _7648_/D vssd2 vssd2 vccd2 vccd2 _7648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_158 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7579_ _7590_/A vssd2 vssd2 vccd2 vccd2 _7579_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_22_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_34_169 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_30_331 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6639__A2 _6040_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5847__B1 _6157_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_30_386 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5362__C _5498_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7049__C1 _7143_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5311__A2 _5528_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5081__D _5468_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5075__A1 _5328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5075__B2 _5145_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4275__A _4898_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_106_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_15_16 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_57_239 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_38_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_108_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_53_445 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6878__A2 _7099_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_111_517 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_504 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7055__A2 _7181_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6950_ _6950_/A _6950_/B vssd2 vssd2 vccd2 vccd2 _6952_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_88_353 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_15_8 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5901_ _7846_/Q _5780_/X _5897_/X _5900_/X _5745_/C vssd2 vssd2 vccd2 vccd2 _5901_/Y
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_0_88_386 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6881_ _6881_/A _6919_/A _6881_/C vssd2 vssd2 vccd2 vccd2 _6919_/B sky130_fd_sc_hd__nand3_1
X_5832_ _7842_/Q _5588_/Y _6017_/B _7844_/Q vssd2 vssd2 vccd2 vccd2 _5832_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_48_228 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_8_336 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5763_ _5769_/B _5763_/B _7871_/Q vssd2 vssd2 vccd2 vccd2 _5764_/C sky130_fd_sc_hd__and3b_1
X_4714_ _4714_/A _4714_/B vssd2 vssd2 vccd2 vccd2 _4717_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__4632__B _5276_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7502_ _7565_/A vssd2 vssd2 vccd2 vccd2 _7502_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_44_456 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5694_ _5694_/A _5694_/B _5694_/C _5694_/D vssd2 vssd2 vccd2 vccd2 _5694_/X sky130_fd_sc_hd__or4_2
XFILLER_0_114_333 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_112_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_71_264 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4645_ _4810_/A _5406_/A _4590_/X _4592_/B vssd2 vssd2 vccd2 vccd2 _4654_/A sky130_fd_sc_hd__o31a_1
X_7433_ hold169/X _7685_/Q _7451_/S vssd2 vssd2 vccd2 vccd2 _7433_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7435__S _7451_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_114_377 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4576_ _4729_/A _5099_/A _5030_/B vssd2 vssd2 vccd2 vccd2 _4581_/A sky130_fd_sc_hd__or3b_2
XANTENNA__5744__A _5781_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7364_ _7440_/A _7364_/B vssd2 vssd2 vccd2 vccd2 _7652_/D sky130_fd_sc_hd__and2_1
Xhold700 _3822_/X vssd2 vssd2 vccd2 vccd2 _3826_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_640 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6315_ _6315_/A _6390_/A vssd2 vssd2 vccd2 vccd2 _6318_/A sky130_fd_sc_hd__nand2_1
X_7295_ _7295_/A _7315_/A vssd2 vssd2 vccd2 vccd2 _7297_/C sky130_fd_sc_hd__nor2_1
X_6246_ _6182_/A _6182_/B _6308_/A vssd2 vssd2 vccd2 vccd2 _6247_/B sky130_fd_sc_hd__a21boi_1
X_6177_ _6177_/A _6177_/B vssd2 vssd2 vccd2 vccd2 _6180_/A sky130_fd_sc_hd__xor2_2
X_5128_ _5128_/A _5128_/B vssd2 vssd2 vccd2 vccd2 _5249_/C sky130_fd_sc_hd__and2_1
XFILLER_0_98_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4807__B _4880_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5059_ _5059_/A _5059_/B vssd2 vssd2 vccd2 vccd2 _5060_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_94_301 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_39_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5919__A _6157_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_109_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_82_507 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_109_149 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_62_220 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5357__C _5357_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_90_584 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_90_562 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5076__D _5076_/D vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_62_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_7_380 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_23_607 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_35_478 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_62_286 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_50_459 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5654__A _7847_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4740__B1 _5406_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_30_194 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6493__B1 _6571_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold82 hold82/A vssd2 vssd2 vccd2 vccd2 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd2 vssd2 vccd2 vccd2 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 hold60/A vssd2 vssd2 vccd2 vccd2 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A vssd2 vssd2 vccd2 vccd2 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_161 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_58_515 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_42_69 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_38_283 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_81_551 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA_2 la_data_in[10] vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_13_139 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4430_ _4427_/X _4429_/X _4022_/B vssd2 vssd2 vccd2 vccd2 _5366_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__5283__B _5404_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_67_11 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6100_ _6094_/B _6281_/B _6282_/A _6100_/D vssd2 vssd2 vccd2 vccd2 _6100_/X sky130_fd_sc_hd__and4b_1
X_4361_ _4420_/A _4361_/B vssd2 vssd2 vccd2 vccd2 _4362_/B sky130_fd_sc_hd__and2_1
X_7080_ _7082_/A vssd2 vssd2 vccd2 vccd2 _7080_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_67_44 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_323 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4292_ _4293_/A _4293_/B vssd2 vssd2 vccd2 vccd2 _4292_/X sky130_fd_sc_hd__and2b_1
X_6031_ _6032_/A _6032_/B vssd2 vssd2 vccd2 vccd2 _6031_/X sky130_fd_sc_hd__or2_1
XTAP_367 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5039__B2 _4962_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_83_87 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_89_673 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XPHY_18 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6933_ _6866_/A _6866_/B _6864_/X vssd2 vssd2 vccd2 vccd2 _6954_/A sky130_fd_sc_hd__a21o_1
X_6864_ _6865_/A _6865_/B vssd2 vssd2 vccd2 vccd2 _6864_/X sky130_fd_sc_hd__and2_1
XFILLER_0_76_378 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5815_ _5816_/A _5816_/B vssd2 vssd2 vccd2 vccd2 _6105_/B sky130_fd_sc_hd__and2_1
XANTENNA__5458__B _5528_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_91_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_6795_ _6795_/A _6795_/B vssd2 vssd2 vccd2 vccd2 _6797_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_592 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5746_ _7845_/Q _6152_/B _6155_/B _5944_/C vssd2 vssd2 vccd2 vccd2 _5760_/A sky130_fd_sc_hd__and4_1
XFILLER_0_32_80 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_44_275 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_44_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5677_ _7875_/Q _7876_/Q vssd2 vssd2 vccd2 vccd2 _5694_/B sky130_fd_sc_hd__or2_4
XFILLER_0_114_141 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7416_ hold212/X _7677_/Q _7418_/S vssd2 vssd2 vccd2 vccd2 _7416_/X sky130_fd_sc_hd__mux2_1
X_4628_ _4814_/A _3971_/Y _4019_/Y _3893_/B _4627_/Y vssd2 vssd2 vccd2 vccd2 _4628_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_32_459 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold530 input17/X vssd2 vssd2 vccd2 vccd2 hold54/A sky130_fd_sc_hd__dlygate4sd3_1
X_4559_ _4500_/A _4500_/B _4501_/Y vssd2 vssd2 vccd2 vccd2 _4573_/A sky130_fd_sc_hd__a21bo_1
Xhold552 la_data_in[44] vssd2 vssd2 vccd2 vccd2 hold67/A sky130_fd_sc_hd__dlygate4sd3_1
X_7347_ hold98/X _7347_/B vssd2 vssd2 vccd2 vccd2 hold99/A sky130_fd_sc_hd__nor2_1
XFILLER_0_13_673 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_40_470 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_40_481 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold563 hold74/X vssd2 vssd2 vccd2 vccd2 _7867_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 hold63/X vssd2 vssd2 vccd2 vccd2 input22/A sky130_fd_sc_hd__dlygate4sd3_1
X_7278_ _7308_/A _7278_/B vssd2 vssd2 vccd2 vccd2 _7283_/A sky130_fd_sc_hd__nand2_1
Xhold585 hold83/X vssd2 vssd2 vccd2 vccd2 input46/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 input43/X vssd2 vssd2 vccd2 vccd2 hold80/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 la_data_in[3] vssd2 vssd2 vccd2 vccd2 hold91/A sky130_fd_sc_hd__dlygate4sd3_1
X_6229_ _6229_/A _6229_/B vssd2 vssd2 vccd2 vccd2 _6233_/A sky130_fd_sc_hd__xnor2_2
XTAP_890 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_79_150 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_79_183 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5450__A1 _4996_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_95_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_94_153 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_82_315 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5202__A1 _5168_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4272__B _5042_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_94_197 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_35_220 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_106_642 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_106_620 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_50_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_2_309 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6662__B _7099_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4463__A _4962_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_53_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3930_ _7762_/Q _4252_/D _4707_/A _3929_/Y vssd2 vssd2 vccd2 vccd2 _3930_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_85_175 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_73_326 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__7194__A1 _7140_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_46_529 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_3861_ _3858_/A _3858_/B _4100_/B vssd2 vssd2 vccd2 vccd2 _3895_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_39_581 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6580_ _6812_/A _6812_/B _7237_/A _7224_/A vssd2 vssd2 vccd2 vccd2 _6582_/B sky130_fd_sc_hd__or4_1
XFILLER_0_73_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5600_ _5594_/X _5599_/X _5588_/Y vssd2 vssd2 vccd2 vccd2 _5600_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_5_103 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_26_231 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_3792_ _4893_/A vssd2 vssd2 vccd2 vccd2 _4814_/A sky130_fd_sc_hd__inv_2
XFILLER_0_54_551 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_26_253 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5531_ _5550_/A _5498_/D _5550_/B _5498_/A vssd2 vssd2 vccd2 vccd2 _5532_/B sky130_fd_sc_hd__o22a_1
XFILLER_0_26_286 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_111_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7201_ _7164_/A _7164_/B _7157_/X vssd2 vssd2 vccd2 vccd2 _7203_/B sky130_fd_sc_hd__o21a_1
X_5462_ _5462_/A _5462_/B vssd2 vssd2 vccd2 vccd2 _5526_/A sky130_fd_sc_hd__or2_1
X_5393_ _5394_/A _5394_/B vssd2 vssd2 vccd2 vccd2 _5393_/X sky130_fd_sc_hd__or2_1
X_4413_ _4413_/A _4413_/B vssd2 vssd2 vccd2 vccd2 _4415_/B sky130_fd_sc_hd__xnor2_2
X_7132_ _7131_/A _7326_/A _7087_/A _7034_/A vssd2 vssd2 vccd2 vccd2 _7133_/B sky130_fd_sc_hd__a31o_1
X_4344_ _4344_/A _4344_/B vssd2 vssd2 vccd2 vccd2 _4345_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_10_643 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7063_ _7064_/A _7064_/B vssd2 vssd2 vccd2 vccd2 _7111_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5741__B _5992_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_94_53 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4275_ _4898_/A _4662_/B _4273_/Y vssd2 vssd2 vccd2 vccd2 _4276_/B sky130_fd_sc_hd__or3b_1
X_6014_ _6074_/A _6194_/C _6130_/C vssd2 vssd2 vccd2 vccd2 _6014_/X sky130_fd_sc_hd__and3_1
XFILLER_0_94_97 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA_fanout274_A _7770_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_96_429 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1319 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_470 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_1308 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6572__B _6572_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_77_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6916_ _6916_/A _6916_/B _6914_/X vssd2 vssd2 vccd2 vccd2 _6916_/X sky130_fd_sc_hd__or3b_1
X_6847_ _6847_/A _6847_/B vssd2 vssd2 vccd2 vccd2 _6847_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_453 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6778_ _6719_/A _6717_/Y _6716_/Y vssd2 vssd2 vccd2 vccd2 _6798_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_9_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_91_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_45_573 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5729_ _7874_/Q _5730_/B vssd2 vssd2 vccd2 vccd2 _5739_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_72_381 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_60_565 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_20_407 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_102_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_60_598 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_60_587 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_20_429 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_102_177 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold360 _7678_/Q vssd2 vssd2 vccd2 vccd2 hold360/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_492 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold371 hold684/X vssd2 vssd2 vccd2 vccd2 _7800_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 hold689/X vssd2 vssd2 vccd2 vccd2 _7777_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _7664_/Q vssd2 vssd2 vccd2 vccd2 hold382/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_87_407 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_114_29 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_95_440 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_68_676 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_67_131 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_95_473 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_55_326 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_55_304 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_23_38 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_55_359 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_106_483 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7479__A2 _7483_/A2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6151__A2 _5816_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4060_ _7764_/Q _4252_/D vssd2 vssd2 vccd2 vccd2 _4060_/Y sky130_fd_sc_hd__nand2_1
X_4962_ _4962_/A _5164_/A _5406_/A _5164_/B vssd2 vssd2 vccd2 vccd2 _5033_/A sky130_fd_sc_hd__or4_2
X_7750_ _7750_/CLK _7750_/D _7509_/Y vssd2 vssd2 vccd2 vccd2 _7750_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_484 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6701_ _6402_/A _7197_/B _6700_/X vssd2 vssd2 vccd2 vccd2 _6754_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_74_602 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_46_304 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4893_ _4893_/A _4893_/B vssd2 vssd2 vccd2 vccd2 _5550_/B sky130_fd_sc_hd__nand2_8
XANTENNA__3976__A1 _4454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3976__B2 _4328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3913_ _7789_/Q _3913_/B vssd2 vssd2 vccd2 vccd2 _3913_/Y sky130_fd_sc_hd__xnor2_2
X_7681_ _7795_/CLK _7681_/D vssd2 vssd2 vccd2 vccd2 _7681_/Q sky130_fd_sc_hd__dfxtp_1
X_6632_ _6576_/A _6576_/C _6576_/B vssd2 vssd2 vccd2 vccd2 _6648_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_58_197 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_6_401 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3844_ _7798_/Q _3844_/B vssd2 vssd2 vccd2 vccd2 _4267_/D sky130_fd_sc_hd__xor2_4
XANTENNA__6914__A1 _6855_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5717__A2 _5992_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_27_551 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6563_ _6563_/A _6563_/B vssd2 vssd2 vccd2 vccd2 _6564_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_223 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6494_ _6571_/A _6571_/C vssd2 vssd2 vccd2 vccd2 _6496_/B sky130_fd_sc_hd__nand2_1
X_5514_ _5515_/A _5515_/B _5515_/C vssd2 vssd2 vccd2 vccd2 _5516_/A sky130_fd_sc_hd__a21oi_1
X_5445_ _5445_/A _5445_/B vssd2 vssd2 vccd2 vccd2 _5445_/X sky130_fd_sc_hd__and2_1
XFILLER_0_14_267 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_112_475 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__7443__S _7451_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4153__A1 _4809_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7115_ _7168_/A _7114_/Y _7047_/A _7197_/B vssd2 vssd2 vccd2 vccd2 _7117_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_10_462 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_1_172 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5376_ _5377_/A _5377_/B vssd2 vssd2 vccd2 vccd2 _5421_/A sky130_fd_sc_hd__nand2_1
X_4327_ _7772_/Q _4075_/B _4325_/X _3827_/Y _4326_/X vssd2 vssd2 vccd2 vccd2 _4327_/X
+ sky130_fd_sc_hd__a221o_2
X_7046_ _7046_/A _7046_/B vssd2 vssd2 vccd2 vccd2 _7048_/A sky130_fd_sc_hd__nand2_1
Xfanout169 _6705_/B vssd2 vssd2 vccd2 vccd2 _6855_/A sky130_fd_sc_hd__clkbuf_8
X_4258_ _4598_/A _4711_/A vssd2 vssd2 vccd2 vccd2 _4260_/C sky130_fd_sc_hd__nor2_1
X_4189_ _4189_/A _4189_/B _4189_/C _4189_/D vssd2 vssd2 vccd2 vccd2 _4190_/A sky130_fd_sc_hd__and4_1
XTAP_1105 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_443 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_64_123 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7879_ _7886_/CLK _7879_/D _7638_/Y vssd2 vssd2 vccd2 vccd2 _7879_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_107_225 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_80_605 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_64_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_64_156 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_521 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_598 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7353__S _7383_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5662__A _6093_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold190 _7431_/X vssd2 vssd2 vccd2 vccd2 _7432_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_237 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4725__B _5315_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_34_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_34_48 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_95_281 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_83_465 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_71_605 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4741__A _4962_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_55_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_113_217 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6668__A _6668_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_67 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5230_ _5231_/A _5231_/B vssd2 vssd2 vccd2 vccd2 _5275_/A sky130_fd_sc_hd__nand2_1
X_5161_ _5162_/A _5162_/B _5162_/C vssd2 vssd2 vccd2 vccd2 _5163_/A sky130_fd_sc_hd__a21o_1
X_5092_ _5090_/X _5092_/B vssd2 vssd2 vccd2 vccd2 _5093_/B sky130_fd_sc_hd__and2b_2
X_4112_ _4110_/Y _4111_/X _4148_/C vssd2 vssd2 vccd2 vccd2 _4112_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_75_77 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5635__A1 _5645_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4043_ _4025_/X _4040_/X _4042_/X _4033_/C vssd2 vssd2 vccd2 vccd2 _4044_/B sky130_fd_sc_hd__o31ai_4
XFILLER_0_59_440 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5994_ _5991_/X _5993_/X _5781_/B vssd2 vssd2 vccd2 vccd2 _5994_/X sky130_fd_sc_hd__o21a_2
X_7802_ _7802_/CLK _7802_/D _7561_/Y vssd2 vssd2 vccd2 vccd2 _7802_/Q sky130_fd_sc_hd__dfrtp_2
X_4945_ _4946_/B _4946_/A vssd2 vssd2 vccd2 vccd2 _4945_/Y sky130_fd_sc_hd__nand2b_1
X_7733_ _7739_/CLK _7733_/D _7492_/Y vssd2 vssd2 vccd2 vccd2 _7733_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_421 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_74_410 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_59_484 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_46_123 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_19_337 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4876_ _4876_/A _4876_/B vssd2 vssd2 vccd2 vccd2 _4877_/B sky130_fd_sc_hd__xnor2_2
X_7664_ _7776_/CLK _7664_/D vssd2 vssd2 vccd2 vccd2 _7664_/Q sky130_fd_sc_hd__dfxtp_1
X_7595_ _7597_/A vssd2 vssd2 vccd2 vccd2 _7595_/Y sky130_fd_sc_hd__inv_2
X_6615_ _6615_/A _6615_/B vssd2 vssd2 vccd2 vccd2 _6615_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_61_126 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3827_ _4809_/B _4893_/B vssd2 vssd2 vccd2 vccd2 _3827_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_27_370 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6546_ _6707_/A _7253_/A _6547_/A vssd2 vssd2 vccd2 vccd2 _6546_/X sky130_fd_sc_hd__or3_1
XFILLER_0_61_159 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XANTENNA__5571__B1 _5548_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_42_373 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6477_ _6542_/A _6477_/B vssd2 vssd2 vccd2 vccd2 _6488_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4126__A1 _4268_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_100_434 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4126__B2 _7766_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5428_ _5363_/A _5365_/B _5363_/B vssd2 vssd2 vccd2 vccd2 _5430_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_100_456 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6728__D _7237_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5359_ _5454_/A _5359_/B vssd2 vssd2 vccd2 vccd2 _7749_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__4098__A _4898_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_100_489 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7029_ _7029_/A _7029_/B vssd2 vssd2 vccd2 vccd2 _7031_/C sky130_fd_sc_hd__and2_1
XFILLER_0_69_215 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_77_292 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_92_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__4561__A _4898_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_108_567 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4280__B _4863_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4711__D _5099_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_18_381 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_20_39 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_21_513 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_110_209 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_60_192 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_261 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5314__B1 _5468_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_708 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4736__A _4736_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_45_47 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_88_513 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_75_218 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6042__A1 _6039_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_0_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6593__A2 _7099_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_56_421 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6670__B _6670_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_1491 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _4730_/A _4730_/B vssd2 vssd2 vccd2 vccd2 _4732_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_424 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4661_ _4662_/B _5099_/A _5315_/B _4807_/A vssd2 vssd2 vccd2 vccd2 _4663_/A sky130_fd_sc_hd__o22ai_1
XFILLER_0_43_104 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_71_468 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6400_ _6396_/Y _6397_/Y _6398_/Y _5653_/C vssd2 vssd2 vccd2 vccd2 _7138_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_43_159 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_9_47 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7380_ _7452_/A _7380_/B vssd2 vssd2 vccd2 vccd2 _7660_/D sky130_fd_sc_hd__and2_1
X_6331_ _6331_/A _6331_/B vssd2 vssd2 vccd2 vccd2 _6332_/B sky130_fd_sc_hd__nor2_1
X_4592_ _4590_/X _4592_/B vssd2 vssd2 vccd2 vccd2 _4593_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_12_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_362 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_24_373 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6262_ _6381_/A _6262_/B vssd2 vssd2 vccd2 vccd2 _6303_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4108__A1 _4809_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_86_65 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5213_ _5213_/A _5213_/B vssd2 vssd2 vccd2 vccd2 _5216_/A sky130_fd_sc_hd__xnor2_1
X_6193_ _7849_/Q _7313_/A _6398_/B _7850_/Q vssd2 vssd2 vccd2 vccd2 _6193_/X sky130_fd_sc_hd__a22o_1
X_5144_ _5145_/A _5145_/B vssd2 vssd2 vccd2 vccd2 _5146_/B sky130_fd_sc_hd__nor2_1
XANTENNA__7022__A _7024_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5075_ _5328_/A _5404_/A _5076_/D _5145_/A vssd2 vssd2 vccd2 vccd2 _5077_/A sky130_fd_sc_hd__o22ai_1
XANTENNA__4646__A _5029_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_79_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4026_ _4252_/B _4252_/D _4214_/C _4164_/C vssd2 vssd2 vccd2 vccd2 _4066_/C sky130_fd_sc_hd__nor4_1
XFILLER_0_29_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6861__A _7047_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_35_80 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_87_590 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__6580__B _6812_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_281 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_59_270 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5977_ _6398_/A _5977_/B vssd2 vssd2 vccd2 vccd2 _5977_/X sky130_fd_sc_hd__and2_1
X_4928_ _4863_/A _5550_/A _4860_/X _4862_/B vssd2 vssd2 vccd2 vccd2 _4930_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_74_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7716_ _7750_/CLK _7716_/D vssd2 vssd2 vccd2 vccd2 _7716_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4595__A1 _4809_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_47_476 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7647_ _7776_/CLK _7647_/D vssd2 vssd2 vccd2 vccd2 _7647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_178 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_34_115 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4859_ _4795_/Y _4804_/B _4804_/A vssd2 vssd2 vccd2 vccd2 _4876_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_34_137 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_105_559 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_105_537 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7578_ _7590_/A vssd2 vssd2 vccd2 vccd2 _7578_/Y sky130_fd_sc_hd__inv_2
X_6529_ _6450_/A _6450_/B _6448_/Y vssd2 vssd2 vccd2 vccd2 _6531_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_30_321 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_42_192 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5847__A1 _6282_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5362__D _5528_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_100_253 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5940__A _7845_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7049__B1 _6281_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5075__A2 _5404_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_97_343 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__7221__B1 _7253_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4586__A1 _4809_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4586__B2 _4268_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_53_402 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_232 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_53_457 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_25_159 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_111_529 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5838__A1 _6283_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_21_387 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XTAP_505 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_79 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__6263__A1 _6138_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7460__B1 _7485_/B1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_88_321 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_72_23 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5900_ _5898_/X _5899_/X _5944_/C vssd2 vssd2 vccd2 vccd2 _5900_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_88_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_48_207 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__6015__B2 _7847_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6015__A1 _7846_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6880_ _7037_/A _7237_/A vssd2 vssd2 vccd2 vccd2 _6881_/C sky130_fd_sc_hd__nor2_1
X_5831_ _5586_/B _5584_/Y _5587_/X _5599_/B _5659_/B vssd2 vssd2 vccd2 vccd2 _6017_/B
+ sky130_fd_sc_hd__o2111a_4
XFILLER_0_91_519 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_8_304 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5762_ _5736_/X _5762_/B _6510_/A _7871_/Q vssd2 vssd2 vccd2 vccd2 _5762_/X sky130_fd_sc_hd__and4b_1
X_4713_ _4896_/A _5276_/A vssd2 vssd2 vccd2 vccd2 _4714_/B sky130_fd_sc_hd__or2_1
XFILLER_0_44_413 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_8_348 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7501_ _7565_/A vssd2 vssd2 vccd2 vccd2 _7501_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_6_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7886_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_44_435 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5693_ _7879_/Q _7880_/Q _7881_/Q _7882_/Q vssd2 vssd2 vccd2 vccd2 _5694_/D sky130_fd_sc_hd__or4_1
XANTENNA__4329__A1 _7767_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4644_ _4581_/A _4581_/B _4579_/Y vssd2 vssd2 vccd2 vccd2 _4655_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__4329__B2 _7766_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_7432_ _7436_/A _7432_/B vssd2 vssd2 vccd2 vccd2 _7684_/D sky130_fd_sc_hd__and2_1
XFILLER_0_25_671 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4575_ _4530_/A _4527_/X _4529_/B vssd2 vssd2 vccd2 vccd2 _4583_/A sky130_fd_sc_hd__o21a_1
X_7363_ hold172/X _7764_/D _7383_/S vssd2 vssd2 vccd2 vccd2 _7363_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_389 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6314_ _6313_/B _6313_/C _6313_/A vssd2 vssd2 vccd2 vccd2 _6390_/A sky130_fd_sc_hd__a21o_1
X_7294_ _7292_/X _7294_/B _7294_/C vssd2 vssd2 vccd2 vccd2 _7315_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_24_192 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6245_ _6245_/A _6245_/B vssd2 vssd2 vccd2 vccd2 _6308_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_387 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_12_365 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XANTENNA__5829__A1 _7847_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4509__C_N _5030_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7451__S _7451_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6176_ _6176_/A _6176_/B vssd2 vssd2 vccd2 vccd2 _6177_/B sky130_fd_sc_hd__xnor2_2
X_5127_ _4993_/A _4993_/B _5067_/A _5067_/B vssd2 vssd2 vccd2 vccd2 _5250_/C sky130_fd_sc_hd__o22a_1
X_5058_ _5059_/A _5059_/B vssd2 vssd2 vccd2 vccd2 _5058_/Y sky130_fd_sc_hd__nor2_1
X_4009_ _4809_/A _4084_/B _3901_/B _4080_/D _4162_/A vssd2 vssd2 vccd2 vccd2 _4009_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_67_516 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_47_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_62_232 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4740__B2 _4807_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6493__A1 _6039_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7361__S _7383_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold50 hold50/A vssd2 vssd2 vccd2 vccd2 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A vssd2 vssd2 vccd2 vccd2 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd2 vssd2 vccd2 vccd2 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd2 vssd2 vccd2 vccd2 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold94 hold94/A vssd2 vssd2 vccd2 vccd2 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_26 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_38_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_81_574 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_26_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_41_405 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7335__C_N _7334_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5228__A2_N _5550_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_3 la_data_in[6] vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5283__C _5406_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_1_502 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4360_ _4360_/A _4360_/B _4360_/C vssd2 vssd2 vccd2 vccd2 _4361_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_111_337 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_324 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4291_ _4291_/A _4291_/B vssd2 vssd2 vccd2 vccd2 _4293_/B sky130_fd_sc_hd__xor2_2
XANTENNA__6484__A1 _6402_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6030_ _6082_/A _6738_/A vssd2 vssd2 vccd2 vccd2 _6032_/B sky130_fd_sc_hd__nand2_1
XTAP_357 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4495__B1 _4782_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_379 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5039__A2 _5468_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_107_51 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_83_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_20_7 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5995__B1 _5781_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_49_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6932_ _6932_/A _6932_/B vssd2 vssd2 vccd2 vccd2 _6956_/A sky130_fd_sc_hd__xnor2_1
XPHY_19 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6863_ _6150_/B _7145_/A _6785_/X _6788_/B vssd2 vssd2 vccd2 vccd2 _6865_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_16_82 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_16_93 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5814_ _5662_/C _5809_/X _5813_/X vssd2 vssd2 vccd2 vccd2 _5816_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_91_305 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_64_519 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_6794_ _6792_/Y _6794_/B vssd2 vssd2 vccd2 vccd2 _6795_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_106_109 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_72_541 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__5755__A _5781_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5745_ _5755_/B _5762_/B _5745_/C vssd2 vssd2 vccd2 vccd2 _5745_/X sky130_fd_sc_hd__and3_1
XFILLER_0_96_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_72_574 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5676_ _7873_/Q _7872_/Q _7871_/Q _7874_/Q vssd2 vssd2 vccd2 vccd2 _5694_/A sky130_fd_sc_hd__or4_4
XFILLER_0_17_468 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_114_153 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7415_ _7450_/A _7415_/B vssd2 vssd2 vccd2 vccd2 _7676_/D sky130_fd_sc_hd__and2_1
X_4627_ _4268_/A _3913_/Y _4252_/D vssd2 vssd2 vccd2 vccd2 _4627_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_384 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
Xhold520 la_data_in[19] vssd2 vssd2 vccd2 vccd2 hold75/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_197 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold553 hold67/X vssd2 vssd2 vccd2 vccd2 input39/A sky130_fd_sc_hd__dlygate4sd3_1
X_4558_ _4558_/A _4558_/B vssd2 vssd2 vccd2 vccd2 _4614_/A sky130_fd_sc_hd__nand2_1
X_7346_ _7346_/A _7346_/B _7346_/C _7346_/D vssd2 vssd2 vccd2 vccd2 _7346_/Y sky130_fd_sc_hd__nor4_1
Xhold531 hold54/X vssd2 vssd2 vccd2 vccd2 _7863_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 input22/X vssd2 vssd2 vccd2 vccd2 hold64/A sky130_fd_sc_hd__dlygate4sd3_1
X_7277_ _7277_/A _7277_/B vssd2 vssd2 vccd2 vccd2 _7278_/B sky130_fd_sc_hd__or2_1
Xhold586 input46/X vssd2 vssd2 vccd2 vccd2 hold84/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 hold91/X vssd2 vssd2 vccd2 vccd2 input34/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 hold80/X vssd2 vssd2 vccd2 vccd2 _7875_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 la_data_in[21] vssd2 vssd2 vccd2 vccd2 hold65/A sky130_fd_sc_hd__dlygate4sd3_1
X_4489_ _4814_/B _4489_/B vssd2 vssd2 vccd2 vccd2 _4489_/X sky130_fd_sc_hd__and2_1
X_6228_ _6228_/A _6228_/B vssd2 vssd2 vccd2 vccd2 _6229_/B sky130_fd_sc_hd__xnor2_2
XTAP_880 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6282_/A _6357_/B _6156_/X _6157_/X _6158_/X vssd2 vssd2 vccd2 vccd2 _6159_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_0_99_405 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XTAP_891 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_94_121 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_94_165 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5202__A2 _5431_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6935__C1 _5992_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5738__B1 _6152_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_90_360 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_63_574 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_23_405 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_90_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_35_276 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_23_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_31_482 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_53_36 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__4463__B _4896_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_46_508 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_85_154 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7194__A2 _7255_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_3860_ _7795_/Q _3860_/B vssd2 vssd2 vccd2 vccd2 _3880_/A sky130_fd_sc_hd__xnor2_2
X_3791_ _7791_/Q vssd2 vssd2 vccd2 vccd2 _3894_/A sky130_fd_sc_hd__inv_2
XPHY_190 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_54_563 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5530_ _5530_/A _5530_/B vssd2 vssd2 vccd2 vccd2 _5532_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_81_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_54_596 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_14_416 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5461_ _5462_/A _5461_/B _5462_/B vssd2 vssd2 vccd2 vccd2 _5463_/B sky130_fd_sc_hd__and3_1
XFILLER_0_78_33 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_7200_ _7242_/A _7200_/B vssd2 vssd2 vccd2 vccd2 _7203_/A sky130_fd_sc_hd__nand2_1
X_4412_ _4412_/A _4412_/B vssd2 vssd2 vccd2 vccd2 _4413_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_55 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5392_ _5392_/A _5392_/B vssd2 vssd2 vccd2 vccd2 _5394_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_41_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_111_167 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7131_ _7131_/A _7131_/B _7131_/C vssd2 vssd2 vccd2 vccd2 _7134_/B sky130_fd_sc_hd__nand3_1
X_4343_ _4044_/A _4044_/B _5042_/B vssd2 vssd2 vccd2 vccd2 _4344_/B sky130_fd_sc_hd__a21oi_2
X_7062_ _7062_/A _7062_/B vssd2 vssd2 vccd2 vccd2 _7064_/B sky130_fd_sc_hd__xnor2_1
X_4274_ _4898_/A _4662_/B _4273_/Y vssd2 vssd2 vccd2 vccd2 _4276_/A sky130_fd_sc_hd__o21bai_2
X_6013_ _6402_/A _6664_/A _5974_/B _5985_/A _5985_/B vssd2 vssd2 vccd2 vccd2 _6026_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_94_65 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6915_ _6916_/A _6916_/B _6914_/X vssd2 vssd2 vccd2 vccd2 _7019_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_11_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6846_ _6847_/A _6847_/B vssd2 vssd2 vccd2 vccd2 _6964_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_443 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_91_113 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6777_ _6707_/A _7291_/B _6901_/A _6776_/X vssd2 vssd2 vccd2 vccd2 _6830_/A sky130_fd_sc_hd__o22ai_4
XFILLER_0_45_552 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5728_ _7873_/Q _7872_/Q _7871_/Q _5735_/B vssd2 vssd2 vccd2 vccd2 _5730_/B sky130_fd_sc_hd__o31a_2
XFILLER_0_17_265 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3989_ _4315_/B _4070_/D _3989_/C _3989_/D vssd2 vssd2 vccd2 vccd2 _3989_/X sky130_fd_sc_hd__and4_1
XFILLER_0_60_533 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5659_ _5659_/A _5659_/B _6019_/C _5811_/B vssd2 vssd2 vccd2 vccd2 _5979_/D sky130_fd_sc_hd__nor4_1
XFILLER_0_60_577 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_13_460 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_20_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7329_ _6588_/B _7197_/B _6669_/X _7313_/A _7315_/A vssd2 vssd2 vccd2 vccd2 _7329_/X
+ sky130_fd_sc_hd__a221o_1
Xhold350 _7483_/X vssd2 vssd2 vccd2 vccd2 _7723_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 _7679_/Q vssd2 vssd2 vccd2 vccd2 hold361/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_189 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
Xhold394 hold687/X vssd2 vssd2 vccd2 vccd2 _7788_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_6 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold383 _7681_/Q vssd2 vssd2 vccd2 vccd2 hold383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 hold683/X vssd2 vssd2 vccd2 vccd2 _7792_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_87_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4564__A _4896_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_67_143 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_67_154 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_55_316 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_28_519 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_82_124 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_36_530 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_63_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_51_566 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_2_107 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_106_495 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_51_577 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_48_25 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6439__A1 _6668_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_48_58 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_31_290 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_wb_clk_i clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2 _7798_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4961_ _5024_/B _4961_/B vssd2 vssd2 vccd2 vccd2 _4978_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_58_121 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_6700_ _6700_/A _6700_/B vssd2 vssd2 vccd2 vccd2 _6700_/X sky130_fd_sc_hd__xor2_1
X_4892_ _4962_/A _5164_/A _5315_/B _5105_/B vssd2 vssd2 vccd2 vccd2 _4958_/A sky130_fd_sc_hd__or4_2
X_3912_ _7789_/Q _3913_/B vssd2 vssd2 vccd2 vccd2 _4068_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_19_519 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7680_ _7795_/CLK _7680_/D vssd2 vssd2 vccd2 vccd2 _7680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_41 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6631_ _6631_/A _6631_/B vssd2 vssd2 vccd2 vccd2 _6650_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_80_67 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_73_135 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_73_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_3843_ _7795_/Q _7796_/Q _7797_/Q _3822_/A _3888_/B vssd2 vssd2 vccd2 vccd2 _3844_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_0_104_85 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_73_146 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6914__A2 _7255_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_6_413 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6562_ _6563_/A _6563_/B vssd2 vssd2 vccd2 vccd2 _6631_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_54_382 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_54_360 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_42_511 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6493_ _6039_/X _6040_/X _6571_/B _5992_/B vssd2 vssd2 vccd2 vccd2 _6496_/A sky130_fd_sc_hd__o211a_1
XFILLER_0_42_533 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5513_ _5541_/B _5513_/B vssd2 vssd2 vccd2 vccd2 _5515_/C sky130_fd_sc_hd__or2_1
XFILLER_0_112_421 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_14_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5444_ _5518_/A vssd2 vssd2 vccd2 vccd2 _5453_/A sky130_fd_sc_hd__inv_2
XFILLER_0_59_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_7114_ _7114_/A _7114_/B _7114_/C vssd2 vssd2 vccd2 vccd2 _7114_/Y sky130_fd_sc_hd__nor3_1
X_5375_ _5325_/A _5550_/B _5373_/Y _5417_/A vssd2 vssd2 vccd2 vccd2 _5377_/B sky130_fd_sc_hd__a2bb2o_1
X_4326_ _4656_/A _4326_/B _4326_/C _4326_/D vssd2 vssd2 vccd2 vccd2 _4326_/X sky130_fd_sc_hd__and4_1
X_7045_ _7045_/A _7140_/A _7253_/A _7253_/B vssd2 vssd2 vccd2 vccd2 _7046_/B sky130_fd_sc_hd__or4_1
XANTENNA__5102__A1 _5220_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4257_ _4250_/X _4251_/X _4256_/X _4214_/C vssd2 vssd2 vccd2 vccd2 _4257_/Y sky130_fd_sc_hd__o31ai_2
X_4188_ _4187_/A _4189_/C _4189_/D vssd2 vssd2 vccd2 vccd2 _4188_/X sky130_fd_sc_hd__a21o_1
XTAP_1117 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_143 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7878_ _7878_/CLK _7878_/D _7637_/Y vssd2 vssd2 vccd2 vccd2 _7878_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_92_411 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6829_ _6829_/A _6829_/B vssd2 vssd2 vccd2 vccd2 _6830_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_64_135 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_64_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_92_477 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_107_237 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_45_393 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_33_555 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_566 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_103_476 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_20_227 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xhold180 input93/X vssd2 vssd2 vccd2 vccd2 hold180/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold191 hold359/X vssd2 vssd2 vccd2 vccd2 _7760_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_87_249 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_83_400 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_95_293 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_68_485 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_55_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_83_477 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_83_499 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_51_330 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_36_382 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_51_352 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clkbuf_leaf_0_wb_clk_i/A vssd2 vssd2 vccd2 vccd2
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_449 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__6668__B _7294_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_59_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
X_5160_ _5160_/A _5160_/B vssd2 vssd2 vccd2 vccd2 _5162_/C sky130_fd_sc_hd__xor2_1
X_5091_ _5091_/A _5091_/B _5089_/Y vssd2 vssd2 vccd2 vccd2 _5092_/B sky130_fd_sc_hd__or3b_1
X_4111_ _4149_/A _4458_/D _4144_/C _4144_/D vssd2 vssd2 vccd2 vccd2 _4111_/X sky130_fd_sc_hd__or4_1
X_4042_ _4268_/A _3943_/X _4018_/A _4025_/D _4041_/X vssd2 vssd2 vccd2 vccd2 _4042_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_91_55 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7801_ _7802_/CLK _7801_/D _7560_/Y vssd2 vssd2 vccd2 vccd2 _7801_/Q sky130_fd_sc_hd__dfrtp_4
X_5993_ _6093_/A _5769_/X _5785_/X _6282_/A _5992_/X vssd2 vssd2 vccd2 vccd2 _5993_/X
+ sky130_fd_sc_hd__a221o_4
X_4944_ _5145_/A _5276_/A _4865_/X _4867_/B vssd2 vssd2 vccd2 vccd2 _4946_/B sky130_fd_sc_hd__o31a_1
X_7732_ _7739_/CLK _7732_/D _7491_/Y vssd2 vssd2 vccd2 vccd2 _7732_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_305 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_59_496 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_46_102 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4071__A1 _4454_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4875_ _4876_/B _4876_/A vssd2 vssd2 vccd2 vccd2 _4875_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_74_455 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_62_617 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_46_135 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7663_ _7793_/CLK _7663_/D vssd2 vssd2 vccd2 vccd2 _7663_/Q sky130_fd_sc_hd__dfxtp_1
X_7594_ _7597_/A vssd2 vssd2 vccd2 vccd2 _7594_/Y sky130_fd_sc_hd__inv_2
X_6614_ _6537_/A _6456_/Y _6537_/B vssd2 vssd2 vccd2 vccd2 _6765_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_105 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_6_232 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_3826_ _3826_/A _3826_/B _3888_/B vssd2 vssd2 vccd2 vccd2 _4006_/B sky130_fd_sc_hd__nor3b_4
X_6545_ _6707_/A _7253_/A vssd2 vssd2 vccd2 vccd2 _6547_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_42_330 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_15_544 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_27_393 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_40_81 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_42_363 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_112_251 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6476_ _6402_/A _7222_/A _7222_/C _5819_/B vssd2 vssd2 vccd2 vccd2 _6477_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_30_525 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XANTENNA__4379__A _4708_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5427_ _5427_/A _5427_/B vssd2 vssd2 vccd2 vccd2 _5433_/A sky130_fd_sc_hd__xnor2_1
X_5358_ _5455_/A _5454_/B vssd2 vssd2 vccd2 vccd2 _5359_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4098__B _4807_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4309_ _5455_/A _4309_/B vssd2 vssd2 vccd2 vccd2 _4362_/A sky130_fd_sc_hd__nand2_1
X_7028_ _6903_/X _6965_/X _6966_/X vssd2 vssd2 vccd2 vccd2 _7029_/B sky130_fd_sc_hd__a21oi_2
X_5289_ _5289_/A _5289_/B vssd2 vssd2 vccd2 vccd2 _5292_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_97_558 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_97_547 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_37_113 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__4561__B _5142_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_65_488 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_53_617 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_18_360 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_37_179 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_80_469 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_80_447 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_20_29 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_33_341 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_0_419 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_21_525 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_21_547 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_103_273 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5314__A1 _5315_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5314__B2 _5404_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_709 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4736__B _5374_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_45_15 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6042__A2 _6040_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_56_411 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_1492 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4660_ _4810_/A _5468_/A vssd2 vssd2 vccd2 vccd2 _4664_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_56_477 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_9_26 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_114_505 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_43_127 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6330_ _6402_/A _6404_/D _6330_/C vssd2 vssd2 vccd2 vccd2 _6331_/B sky130_fd_sc_hd__and3_1
X_4591_ _4962_/A _4662_/B _5042_/B _5222_/A vssd2 vssd2 vccd2 vccd2 _4592_/B sky130_fd_sc_hd__or4_1
XFILLER_0_24_385 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_6261_ _6261_/A _6261_/B _6261_/C vssd2 vssd2 vccd2 vccd2 _6262_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_3_279 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5212_ _5276_/A _5406_/A vssd2 vssd2 vccd2 vccd2 _5213_/B sky130_fd_sc_hd__nor2_1
X_6192_ _6397_/A _6016_/B _6071_/B _6017_/B _6074_/A vssd2 vssd2 vccd2 vccd2 _6192_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_86_77 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_5143_ _5143_/A _5201_/A vssd2 vssd2 vccd2 vccd2 _5146_/A sky130_fd_sc_hd__nand2_1
X_5074_ _5022_/A _5020_/Y _5019_/Y vssd2 vssd2 vccd2 vccd2 _5093_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__4646__B _5222_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4816__B1 _5528_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7022__B _7024_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_4025_ _4018_/A _3965_/A _4025_/C _4025_/D vssd2 vssd2 vccd2 vccd2 _4025_/X sky130_fd_sc_hd__and4bb_1
XFILLER_0_79_558 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__7449__S _7451_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6861__B _7145_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6580__C _7237_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4662__A _4807_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5976_ _7845_/Q _7313_/A _6398_/B _7846_/Q vssd2 vssd2 vccd2 vccd2 _5976_/X sky130_fd_sc_hd__a22o_1
X_4927_ _4877_/A _4877_/B _4875_/X vssd2 vssd2 vccd2 vccd2 _4930_/A sky130_fd_sc_hd__a21oi_1
X_7715_ _7750_/CLK _7715_/D vssd2 vssd2 vccd2 vccd2 _7715_/Q sky130_fd_sc_hd__dfxtp_1
X_4858_ _4787_/A _4787_/B _4788_/Y vssd2 vssd2 vccd2 vccd2 _4877_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_62_425 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7646_ _7776_/CLK _7646_/D vssd2 vssd2 vccd2 vccd2 _7646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_505 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_3809_ _3888_/B _7801_/Q vssd2 vssd2 vccd2 vccd2 _3811_/C sky130_fd_sc_hd__and2_1
XFILLER_0_34_127 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7577_ _7590_/A vssd2 vssd2 vccd2 vccd2 _7577_/Y sky130_fd_sc_hd__inv_2
X_4789_ _4789_/A _4789_/B vssd2 vssd2 vccd2 vccd2 _4791_/B sky130_fd_sc_hd__xnor2_4
X_6528_ _6528_/A _6528_/B vssd2 vssd2 vccd2 vccd2 _6531_/A sky130_fd_sc_hd__xnor2_2
X_6459_ _6390_/B _6387_/Y _6389_/B vssd2 vssd2 vccd2 vccd2 _6461_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_100_221 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5847__A2 _5992_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_100_265 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__7221__A1 _7291_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7359__S _7383_/S vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7221__B2 _7253_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4035__A1 _7764_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_38_400 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_108_321 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_53_414 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_38_477 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_108_365 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_80_266 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_34_661 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_34_672 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_40_108 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_33_193 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XTAP_506 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4747__A _4747_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__6263__A2 _6973_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4274__A1 _4898_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_76_517 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_76_506 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_72_68 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_76_539 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5830_ _5599_/B _5653_/C _5829_/X _6474_/A _7843_/Q vssd2 vssd2 vccd2 vccd2 _5830_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_400 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_91_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_56_241 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5774__A1 _7845_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5774__B2 _7847_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5761_ _5717_/X _5737_/Y _5745_/X _5736_/X _5760_/X vssd2 vssd2 vccd2 vccd2 _5761_/X
+ sky130_fd_sc_hd__a221o_1
X_4712_ _4712_/A _4712_/B vssd2 vssd2 vccd2 vccd2 _4714_/A sky130_fd_sc_hd__nand2_1
X_7500_ _7561_/A vssd2 vssd2 vccd2 vccd2 _7500_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_112_41 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_5692_ _5691_/A _5691_/B _5937_/B vssd2 vssd2 vccd2 vccd2 _6152_/C sky130_fd_sc_hd__a21oi_4
XFILLER_0_16_138 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7431_ hold172/X _7796_/D _7451_/S vssd2 vssd2 vccd2 vccd2 _7431_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_112_85 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
X_4643_ _4643_/A _4643_/B vssd2 vssd2 vccd2 vccd2 _4677_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_50 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_4574_ _4514_/A _4514_/B _4512_/Y vssd2 vssd2 vccd2 vccd2 _4584_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_12_300 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7362_ _7440_/A _7362_/B vssd2 vssd2 vccd2 vccd2 _7651_/D sky130_fd_sc_hd__and2_1
XFILLER_0_31_119 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_6313_ _6313_/A _6313_/B _6313_/C vssd2 vssd2 vccd2 vccd2 _6315_/A sky130_fd_sc_hd__nand3_1
X_7293_ _7253_/C _7255_/B _7292_/X vssd2 vssd2 vccd2 vccd2 _7295_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_12_333 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6244_ _6245_/A _6245_/B vssd2 vssd2 vccd2 vccd2 _6387_/A sky130_fd_sc_hd__nor2_1
X_6175_ _6176_/B _6176_/A vssd2 vssd2 vccd2 vccd2 _6175_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_41_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_5126_ _5126_/A _5126_/B vssd2 vssd2 vccd2 vccd2 _5250_/B sky130_fd_sc_hd__xnor2_4
X_5057_ _4982_/A _4982_/B _4980_/X vssd2 vssd2 vccd2 vccd2 _5059_/B sky130_fd_sc_hd__a21oi_4
X_4008_ _4519_/C _4267_/C _4267_/D vssd2 vssd2 vccd2 vccd2 _4200_/B sky130_fd_sc_hd__and3_1
XANTENNA__4265__B2 _7767_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4265__A1 _4328_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4397__A_N _4896_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_94_369 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_5959_ _5958_/B _5958_/C _5958_/A vssd2 vssd2 vccd2 vccd2 _5960_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_572 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_75_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_35_414 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_90_542 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_105_335 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_7629_ _7629_/A vssd2 vssd2 vccd2 vccd2 _7629_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_35_458 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_50_417 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XANTENNA__4740__A2 _4965_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_30_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_30_152 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6493__A2 _6040_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold40 hold40/A vssd2 vssd2 vccd2 vccd2 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd2 vssd2 vccd2 vccd2 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd2 vssd2 vccd2 vccd2 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_39 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
Xhold73 hold73/A vssd2 vssd2 vccd2 vccd2 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd2 vssd2 vccd2 vccd2 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd2 vssd2 vccd2 vccd2 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5756__A1 _6158_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__5756__B2 _6283_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_81_531 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_108_195 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_81_586 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_53_277 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_41_417 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_0_111_305 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__5283__D _5498_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA_4 la_data_in[9] vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_34_491 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_111_349 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_67_57 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
X_4290_ _4291_/A _4291_/B vssd2 vssd2 vccd2 vccd2 _4351_/A sky130_fd_sc_hd__nand2_1
XTAP_314 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6484__A2 _7145_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4495__A1 _4896_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_358 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4495__B2 _4704_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XTAP_369 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_152 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_88_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5995__A1 _5991_/X vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_6931_ _6932_/A _6932_/B vssd2 vssd2 vccd2 vccd2 _7007_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_7 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_16_61 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_6862_ _6862_/A _6862_/B vssd2 vssd2 vccd2 vccd2 _6865_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_64_509 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5813_ _7844_/Q _5812_/C _5810_/X _5812_/X _5663_/X vssd2 vssd2 vccd2 vccd2 _5813_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_91_317 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_57_572 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_6793_ _6793_/A _6793_/B vssd2 vssd2 vccd2 vccd2 _6794_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4940__A _5210_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
X_5744_ _5781_/B _5744_/B _5755_/C _5936_/B vssd2 vssd2 vccd2 vccd2 _5745_/C sky130_fd_sc_hd__nor4b_4
X_5675_ _6436_/A vssd2 vssd2 vccd2 vccd2 _6105_/A sky130_fd_sc_hd__inv_2
XFILLER_0_72_553 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_89_3 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_72_586 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_4626_ _4584_/A _4584_/B _4582_/Y vssd2 vssd2 vccd2 vccd2 _4641_/A sky130_fd_sc_hd__a21o_1
X_7414_ hold194/X _7676_/Q _7418_/S vssd2 vssd2 vccd2 vccd2 _7414_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_165 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
Xhold510 input42/X vssd2 vssd2 vccd2 vccd2 hold40/A sky130_fd_sc_hd__dlygate4sd3_1
X_7345_ _7345_/A _7345_/B _7345_/C _7345_/D vssd2 vssd2 vccd2 vccd2 _7346_/D sky130_fd_sc_hd__or4_1
Xhold554 input39/X vssd2 vssd2 vccd2 vccd2 hold68/A sky130_fd_sc_hd__dlygate4sd3_1
X_4557_ _5455_/A _4557_/B vssd2 vssd2 vccd2 vccd2 _4622_/A sky130_fd_sc_hd__nand2_1
Xmax_cap240 _3967_/C vssd2 vssd2 vccd2 vccd2 _4036_/B sky130_fd_sc_hd__buf_1
Xhold521 hold75/X vssd2 vssd2 vccd2 vccd2 input11/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 la_data_in[25] vssd2 vssd2 vccd2 vccd2 hold57/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 hold64/X vssd2 vssd2 vccd2 vccd2 _7868_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_450 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_7276_ _7277_/A _7277_/B vssd2 vssd2 vccd2 vccd2 _7308_/A sky130_fd_sc_hd__nand2_1
Xhold576 la_data_in[6] vssd2 vssd2 vccd2 vccd2 hold81/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 hold84/X vssd2 vssd2 vccd2 vccd2 _7878_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 hold65/X vssd2 vssd2 vccd2 vccd2 input14/A sky130_fd_sc_hd__dlygate4sd3_1
X_4488_ _7771_/Q _4707_/A _3928_/X _7772_/Q vssd2 vssd2 vccd2 vccd2 _4489_/B sky130_fd_sc_hd__a22o_1
X_6227_ _6590_/A _6228_/A _7197_/A vssd2 vssd2 vccd2 vccd2 _6227_/X sky130_fd_sc_hd__and3_1
XANTENNA__4387__A _4810_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
Xhold598 input34/X vssd2 vssd2 vccd2 vccd2 hold92/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_870 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6158_/A _6283_/B _6587_/B vssd2 vssd2 vccd2 vccd2 _6158_/X sky130_fd_sc_hd__and3_1
XFILLER_0_99_428 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XTAP_892 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _5110_/B _5110_/A vssd2 vssd2 vccd2 vccd2 _5109_/X sky130_fd_sc_hd__and2b_1
XTAP_881 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ _6812_/A _6783_/A _6812_/B _6855_/A vssd2 vssd2 vccd2 vccd2 _6090_/B sky130_fd_sc_hd__or4_1
XFILLER_0_94_133 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XANTENNA__5011__A _5011_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_94_177 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XANTENNA__6935__B1 _7222_/C vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__4850__A _5455_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_23_417 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_50_258 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_16_491 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__4174__B1 _5042_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__3921__B1 _4050_/B vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XANTENNA__7401__A _7440_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_58_325 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_0_58_314 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_58_303 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_53_48 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__6017__A _6157_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_85_111 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_0_73_317 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XANTENNA__5856__A _6283_/A vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_39_561 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_191 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_180 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_54_586 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
X_5460_ _5461_/B _5462_/B vssd2 vssd2 vccd2 vccd2 _5463_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_112_625 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_4411_ _4412_/A _4412_/B vssd2 vssd2 vccd2 vccd2 _4411_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_111_113 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_78_67 vssd2 vssd2 vccd2 vccd2 sky130_ef_sc_hd__decap_12
XFILLER_0_78_45 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
X_5391_ _5344_/A _5343_/Y _5338_/X vssd2 vssd2 vccd2 vccd2 _5392_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__5901__A1 _7846_/Q vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__diode_2
XFILLER_0_22_450 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
X_7130_ _7211_/C _7130_/B vssd2 vssd2 vccd2 vccd2 _7134_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_78_89 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
X_4342_ _5029_/A _4896_/A vssd2 vssd2 vccd2 vccd2 _4344_/A sky130_fd_sc_hd__nor2_2
X_7061_ _7062_/B _7062_/A vssd2 vssd2 vccd2 vccd2 _7114_/B sky130_fd_sc_hd__and2b_1
X_4273_ _4962_/A _4896_/A vssd2 vssd2 vccd2 vccd2 _4273_/Y sky130_fd_sc_hd__nor2_1
X_6012_ _6008_/A _6007_/B _6005_/X vssd2 vssd2 vccd2 vccd2 _6057_/A sky130_fd_sc_hd__a21o_1
.ends

