// This is the unpowered netlist.
module user_proj_example (wb_clk_i,
    io_in,
    io_oeb,
    io_out);
 input wb_clk_i;
 input [6:0] io_in;
 output [6:0] io_oeb;
 output [6:0] io_out;

 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf_wb_clk_i;
 wire net1;
 wire net2;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net5;
 wire net6;
 wire net7;
 wire \top_module_inst.nbit_counter_inst.count0[0] ;
 wire \top_module_inst.nbit_counter_inst.count0[1] ;
 wire \top_module_inst.nbit_counter_inst.count0[2] ;
 wire \top_module_inst.nbit_counter_inst.count0[3] ;
 wire \top_module_inst.nbit_counter_inst.count0[4] ;
 wire \top_module_inst.nbit_counter_inst.count1[0] ;
 wire \top_module_inst.nbit_counter_inst.count1[1] ;
 wire \top_module_inst.nbit_counter_inst.count1[2] ;
 wire \top_module_inst.nbit_counter_inst.count1[3] ;
 wire \top_module_inst.nbit_counter_inst.count1[4] ;
 wire \top_module_inst.nbit_counter_inst.fl ;

 sky130_fd_sc_hd__diode_2 ANTENNA__082__A3 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__083__A_N (.DIODE(_032_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold18_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_output7_A (.DIODE(net7));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_0_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_0_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_100_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_102_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_102_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_105_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_108_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_108_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_109_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_10_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_10_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_110_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_110_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_111_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_111_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_111_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_111_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_111_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_111_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_111_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_111_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_111_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_111_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_111_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_111_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_111_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_111_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_111_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_111_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1034 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_112_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_981 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_1036 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_1044 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_114_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_115_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_1024 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_116_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1033 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_953 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_117_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_117_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_118_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_981 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_118_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1013 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1024 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_119_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_119_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_11_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1047 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120_985 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_120_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1017 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_975 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_122_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_122_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_122_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_122_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_122_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_122_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_122_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_122_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_122_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_122_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_122_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_122_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_122_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_122_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_122_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_122_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_122_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_122_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_123_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_123_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_123_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_123_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_123_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_123_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_123_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_123_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_123_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_123_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_123_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_123_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_123_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_123_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_123_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_123_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_123_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_1017 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_125_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_125_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_126_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_126_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_127_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_128_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_130_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_132_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_133_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_134_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_134_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_136_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_138_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_139_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_13_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_13_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_140_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_142_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_142_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_143_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_143_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_144_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_145_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_146_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_147_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_147_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_148_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_149_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_149_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_14_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_150_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_150_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_153_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_153_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_154_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_154_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_155_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_156_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_157_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_157_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_158_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_15_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_160_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_161_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_161_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_162_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_162_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_163_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_1033 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_164_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_164_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_165_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_165_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_166_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_168_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_170_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_170_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_171_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_172_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_173_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_173_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_174_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_174_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_17_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_17_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_18_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_18_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_20_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_21_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_21_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_22_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_23_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_25_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_25_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_26_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_26_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_27_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_27_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_28_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_28_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_29_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_2_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_2_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_30_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_30_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_32_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_33_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_33_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_34_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_35_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_35_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_36_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_37_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_38_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_3_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_3_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_40_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_41_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_42_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_43_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_43_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_44_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_44_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_45_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_48_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_49_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_4_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_50_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_51_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_51_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_1033 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_53_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_54_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_55_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_57_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_58_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_58_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_59_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_59_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_5_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_5_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_60_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_60_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_62_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_62_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_63_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_63_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_65_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_65_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_66_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_66_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_67_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_67_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_6_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_6_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_70_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_70_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_71_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_71_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_72_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_73_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_73_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_74_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_75_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_76_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_78_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_79_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_79_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_81_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_81_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_82_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_83_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_84_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_86_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_87_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_87_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_88_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_89_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_89_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_90_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_90_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_92_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_92_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_93_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_93_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_95_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_95_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_97_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_98_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_98_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_9_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_9_993 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _076_ (.A(net35),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _077_ (.A(\top_module_inst.nbit_counter_inst.count1[1] ),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _078_ (.A(\top_module_inst.nbit_counter_inst.count0[1] ),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _079_ (.A(net40),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _080_ (.A(net25),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _081_ (.A(net6),
    .Y(_001_));
 sky130_fd_sc_hd__o31a_1 _082_ (.A1(net3),
    .A2(net2),
    .A3(net1),
    .B1(net4),
    .X(_032_));
 sky130_fd_sc_hd__and2b_2 _083_ (.A_N(_032_),
    .B(net5),
    .X(_033_));
 sky130_fd_sc_hd__inv_2 _084_ (.A(_033_),
    .Y(_034_));
 sky130_fd_sc_hd__and2b_1 _085_ (.A_N(net23),
    .B(net21),
    .X(_035_));
 sky130_fd_sc_hd__and2b_1 _086_ (.A_N(net21),
    .B(net23),
    .X(_036_));
 sky130_fd_sc_hd__nor2_1 _087_ (.A(_035_),
    .B(_036_),
    .Y(_037_));
 sky130_fd_sc_hd__o211a_1 _088_ (.A1(\top_module_inst.nbit_counter_inst.count1[3] ),
    .A2(\top_module_inst.nbit_counter_inst.count0[3] ),
    .B1(\top_module_inst.nbit_counter_inst.count0[2] ),
    .C1(\top_module_inst.nbit_counter_inst.count1[2] ),
    .X(_038_));
 sky130_fd_sc_hd__a211o_1 _089_ (.A1(\top_module_inst.nbit_counter_inst.count1[3] ),
    .A2(\top_module_inst.nbit_counter_inst.count0[3] ),
    .B1(_038_),
    .C1(\top_module_inst.nbit_counter_inst.count1[1] ),
    .X(_039_));
 sky130_fd_sc_hd__xor2_1 _090_ (.A(_037_),
    .B(_039_),
    .X(_040_));
 sky130_fd_sc_hd__nor2_1 _091_ (.A(\top_module_inst.nbit_counter_inst.count1[2] ),
    .B(\top_module_inst.nbit_counter_inst.count0[2] ),
    .Y(_041_));
 sky130_fd_sc_hd__xor2_1 _092_ (.A(\top_module_inst.nbit_counter_inst.count1[2] ),
    .B(\top_module_inst.nbit_counter_inst.count0[2] ),
    .X(_042_));
 sky130_fd_sc_hd__xor2_1 _093_ (.A(net41),
    .B(\top_module_inst.nbit_counter_inst.count0[0] ),
    .X(_043_));
 sky130_fd_sc_hd__nand2b_1 _094_ (.A_N(\top_module_inst.nbit_counter_inst.count1[1] ),
    .B(\top_module_inst.nbit_counter_inst.count0[1] ),
    .Y(_044_));
 sky130_fd_sc_hd__o211a_1 _095_ (.A1(_028_),
    .A2(_042_),
    .B1(net42),
    .C1(_044_),
    .X(_045_));
 sky130_fd_sc_hd__xor2_1 _096_ (.A(net35),
    .B(net30),
    .X(_046_));
 sky130_fd_sc_hd__a2bb2o_1 _097_ (.A1_N(_041_),
    .A2_N(_046_),
    .B1(_042_),
    .B2(_029_),
    .X(_047_));
 sky130_fd_sc_hd__a21o_1 _098_ (.A1(_041_),
    .A2(_046_),
    .B1(_047_),
    .X(_048_));
 sky130_fd_sc_hd__or3b_2 _099_ (.A(_048_),
    .B(_040_),
    .C_N(_045_),
    .X(_049_));
 sky130_fd_sc_hd__a21o_1 _100_ (.A1(_034_),
    .A2(_049_),
    .B1(_031_),
    .X(_050_));
 sky130_fd_sc_hd__nand2_1 _101_ (.A(net37),
    .B(net34),
    .Y(_051_));
 sky130_fd_sc_hd__and3_1 _102_ (.A(net26),
    .B(\top_module_inst.nbit_counter_inst.count1[1] ),
    .C(net34),
    .X(_052_));
 sky130_fd_sc_hd__inv_2 _103_ (.A(_052_),
    .Y(_053_));
 sky130_fd_sc_hd__nand2_1 _104_ (.A(net35),
    .B(_052_),
    .Y(_054_));
 sky130_fd_sc_hd__nor2_1 _105_ (.A(net23),
    .B(_031_),
    .Y(_055_));
 sky130_fd_sc_hd__mux2_1 _106_ (.A0(_055_),
    .A1(net23),
    .S(_054_),
    .X(_056_));
 sky130_fd_sc_hd__a32o_1 _107_ (.A1(_033_),
    .A2(_049_),
    .A3(_056_),
    .B1(_050_),
    .B2(net23),
    .X(_023_));
 sky130_fd_sc_hd__or2_1 _108_ (.A(net35),
    .B(_052_),
    .X(_057_));
 sky130_fd_sc_hd__and3_1 _109_ (.A(net25),
    .B(_033_),
    .C(_049_),
    .X(_058_));
 sky130_fd_sc_hd__a32o_1 _110_ (.A1(_054_),
    .A2(_057_),
    .A3(_058_),
    .B1(_050_),
    .B2(net35),
    .X(_022_));
 sky130_fd_sc_hd__a21o_1 _111_ (.A1(\top_module_inst.nbit_counter_inst.count1[1] ),
    .A2(\top_module_inst.nbit_counter_inst.count1[0] ),
    .B1(net26),
    .X(_059_));
 sky130_fd_sc_hd__a32o_1 _112_ (.A1(_053_),
    .A2(_058_),
    .A3(_059_),
    .B1(_050_),
    .B2(net26),
    .X(_021_));
 sky130_fd_sc_hd__or2_1 _113_ (.A(net37),
    .B(net34),
    .X(_060_));
 sky130_fd_sc_hd__a32o_1 _114_ (.A1(_051_),
    .A2(_058_),
    .A3(_060_),
    .B1(_050_),
    .B2(net37),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _115_ (.A0(_058_),
    .A1(_050_),
    .S(net34),
    .X(_019_));
 sky130_fd_sc_hd__or2_1 _116_ (.A(_031_),
    .B(net43),
    .X(_061_));
 sky130_fd_sc_hd__nand2b_1 _117_ (.A_N(net26),
    .B(net28),
    .Y(_062_));
 sky130_fd_sc_hd__and2b_1 _118_ (.A_N(\top_module_inst.nbit_counter_inst.count0[1] ),
    .B(net37),
    .X(_063_));
 sky130_fd_sc_hd__a311o_1 _119_ (.A1(net34),
    .A2(_030_),
    .A3(_044_),
    .B1(_063_),
    .C1(_042_),
    .X(_064_));
 sky130_fd_sc_hd__a21oi_1 _120_ (.A1(_062_),
    .A2(_064_),
    .B1(_046_),
    .Y(_065_));
 sky130_fd_sc_hd__a21oi_1 _121_ (.A1(_027_),
    .A2(net30),
    .B1(_065_),
    .Y(_066_));
 sky130_fd_sc_hd__o21ba_1 _122_ (.A1(_036_),
    .A2(_066_),
    .B1_N(_035_),
    .X(_067_));
 sky130_fd_sc_hd__mux2_1 _123_ (.A0(_067_),
    .A1(net38),
    .S(_061_),
    .X(_018_));
 sky130_fd_sc_hd__nand2_1 _124_ (.A(net32),
    .B(\top_module_inst.nbit_counter_inst.count0[0] ),
    .Y(_068_));
 sky130_fd_sc_hd__and3_1 _125_ (.A(net28),
    .B(\top_module_inst.nbit_counter_inst.count0[1] ),
    .C(\top_module_inst.nbit_counter_inst.count0[0] ),
    .X(_069_));
 sky130_fd_sc_hd__inv_2 _126_ (.A(_069_),
    .Y(_070_));
 sky130_fd_sc_hd__nand2_1 _127_ (.A(net30),
    .B(_069_),
    .Y(_071_));
 sky130_fd_sc_hd__nor2_1 _128_ (.A(net21),
    .B(_031_),
    .Y(_072_));
 sky130_fd_sc_hd__mux2_1 _129_ (.A0(_072_),
    .A1(net21),
    .S(_071_),
    .X(_073_));
 sky130_fd_sc_hd__a21o_1 _130_ (.A1(_033_),
    .A2(_049_),
    .B1(_031_),
    .X(_074_));
 sky130_fd_sc_hd__a32o_1 _131_ (.A1(_034_),
    .A2(_049_),
    .A3(_073_),
    .B1(_074_),
    .B2(net21),
    .X(_017_));
 sky130_fd_sc_hd__or2_1 _132_ (.A(net30),
    .B(_069_),
    .X(_075_));
 sky130_fd_sc_hd__and3_1 _133_ (.A(net25),
    .B(_034_),
    .C(_049_),
    .X(_024_));
 sky130_fd_sc_hd__a32o_1 _134_ (.A1(_071_),
    .A2(_075_),
    .A3(_024_),
    .B1(_074_),
    .B2(net30),
    .X(_016_));
 sky130_fd_sc_hd__a21o_1 _135_ (.A1(\top_module_inst.nbit_counter_inst.count0[1] ),
    .A2(\top_module_inst.nbit_counter_inst.count0[0] ),
    .B1(net28),
    .X(_025_));
 sky130_fd_sc_hd__a32o_1 _136_ (.A1(_070_),
    .A2(_024_),
    .A3(_025_),
    .B1(_074_),
    .B2(net28),
    .X(_015_));
 sky130_fd_sc_hd__or2_1 _137_ (.A(net32),
    .B(\top_module_inst.nbit_counter_inst.count0[0] ),
    .X(_026_));
 sky130_fd_sc_hd__a32o_1 _138_ (.A1(_068_),
    .A2(_024_),
    .A3(_026_),
    .B1(_074_),
    .B2(net32),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _139_ (.A0(_074_),
    .A1(_024_),
    .S(_030_),
    .X(_013_));
 sky130_fd_sc_hd__o21a_1 _140_ (.A1(net25),
    .A2(_033_),
    .B1(_061_),
    .X(_000_));
 sky130_fd_sc_hd__inv_2 _141_ (.A(net6),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _142_ (.A(net6),
    .Y(_003_));
 sky130_fd_sc_hd__inv_2 _143_ (.A(net6),
    .Y(_004_));
 sky130_fd_sc_hd__inv_2 _144_ (.A(net6),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _145_ (.A(net6),
    .Y(_006_));
 sky130_fd_sc_hd__inv_2 _146_ (.A(net6),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _147_ (.A(net6),
    .Y(_008_));
 sky130_fd_sc_hd__inv_2 _148_ (.A(net6),
    .Y(_009_));
 sky130_fd_sc_hd__inv_2 _149_ (.A(net6),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _150_ (.A(net6),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _151_ (.A(net6),
    .Y(_012_));
 sky130_fd_sc_hd__dfrtp_2 _152_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(_013_),
    .RESET_B(_001_),
    .Q(\top_module_inst.nbit_counter_inst.count0[0] ));
 sky130_fd_sc_hd__dfrtp_2 _153_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(net33),
    .RESET_B(_002_),
    .Q(\top_module_inst.nbit_counter_inst.count0[1] ));
 sky130_fd_sc_hd__dfrtp_2 _154_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(net29),
    .RESET_B(_003_),
    .Q(\top_module_inst.nbit_counter_inst.count0[2] ));
 sky130_fd_sc_hd__dfrtp_1 _155_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(net31),
    .RESET_B(_004_),
    .Q(\top_module_inst.nbit_counter_inst.count0[3] ));
 sky130_fd_sc_hd__dfrtp_1 _156_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(net22),
    .RESET_B(_005_),
    .Q(\top_module_inst.nbit_counter_inst.count0[4] ));
 sky130_fd_sc_hd__dfrtp_2 _157_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(net39),
    .RESET_B(_006_),
    .Q(net7));
 sky130_fd_sc_hd__dfrtp_1 _158_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(_019_),
    .RESET_B(_007_),
    .Q(\top_module_inst.nbit_counter_inst.count1[0] ));
 sky130_fd_sc_hd__dfrtp_2 _159_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(_020_),
    .RESET_B(_008_),
    .Q(\top_module_inst.nbit_counter_inst.count1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _160_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(net27),
    .RESET_B(_009_),
    .Q(\top_module_inst.nbit_counter_inst.count1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _161_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(net36),
    .RESET_B(_010_),
    .Q(\top_module_inst.nbit_counter_inst.count1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _162_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(net24),
    .RESET_B(_011_),
    .Q(\top_module_inst.nbit_counter_inst.count1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _163_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(_000_),
    .RESET_B(_012_),
    .Q(\top_module_inst.nbit_counter_inst.fl ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__buf_1 hold1 (.A(\top_module_inst.nbit_counter_inst.count0[4] ),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 hold10 (.A(\top_module_inst.nbit_counter_inst.count0[3] ),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_016_),
    .X(net31));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\top_module_inst.nbit_counter_inst.count0[1] ),
    .X(net32));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_014_),
    .X(net33));
 sky130_fd_sc_hd__buf_1 hold14 (.A(net45),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 hold15 (.A(\top_module_inst.nbit_counter_inst.count1[3] ),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_022_),
    .X(net36));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold17 (.A(\top_module_inst.nbit_counter_inst.count1[1] ),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net7),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_018_),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_017_),
    .X(net22));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\top_module_inst.nbit_counter_inst.count0[0] ),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\top_module_inst.nbit_counter_inst.count1[0] ),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_043_),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_049_),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\top_module_inst.nbit_counter_inst.fl ),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\top_module_inst.nbit_counter_inst.count1[0] ),
    .X(net45));
 sky130_fd_sc_hd__buf_1 hold3 (.A(\top_module_inst.nbit_counter_inst.count1[4] ),
    .X(net23));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_023_),
    .X(net24));
 sky130_fd_sc_hd__buf_1 hold5 (.A(net44),
    .X(net25));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\top_module_inst.nbit_counter_inst.count1[2] ),
    .X(net26));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_021_),
    .X(net27));
 sky130_fd_sc_hd__buf_1 hold8 (.A(\top_module_inst.nbit_counter_inst.count0[2] ),
    .X(net28));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_015_),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(io_in[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(io_in[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_8 input6 (.A(io_in[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_12 output7 (.A(net7),
    .X(io_out[6]));
 sky130_fd_sc_hd__conb_1 user_proj_example_10 (.LO(net10));
 sky130_fd_sc_hd__conb_1 user_proj_example_11 (.LO(net11));
 sky130_fd_sc_hd__conb_1 user_proj_example_12 (.LO(net12));
 sky130_fd_sc_hd__conb_1 user_proj_example_13 (.LO(net13));
 sky130_fd_sc_hd__conb_1 user_proj_example_14 (.LO(net14));
 sky130_fd_sc_hd__conb_1 user_proj_example_15 (.HI(net15));
 sky130_fd_sc_hd__conb_1 user_proj_example_16 (.HI(net16));
 sky130_fd_sc_hd__conb_1 user_proj_example_17 (.HI(net17));
 sky130_fd_sc_hd__conb_1 user_proj_example_18 (.HI(net18));
 sky130_fd_sc_hd__conb_1 user_proj_example_19 (.HI(net19));
 sky130_fd_sc_hd__conb_1 user_proj_example_20 (.HI(net20));
 sky130_fd_sc_hd__conb_1 user_proj_example_8 (.LO(net8));
 sky130_fd_sc_hd__conb_1 user_proj_example_9 (.LO(net9));
 assign io_oeb[0] = net15;
 assign io_oeb[1] = net16;
 assign io_oeb[2] = net17;
 assign io_oeb[3] = net18;
 assign io_oeb[4] = net19;
 assign io_oeb[5] = net20;
 assign io_oeb[6] = net8;
 assign io_out[0] = net9;
 assign io_out[1] = net10;
 assign io_out[2] = net11;
 assign io_out[3] = net12;
 assign io_out[4] = net13;
 assign io_out[5] = net14;
endmodule

